// Generator : SpinalHDL v1.8.1    git head : 2a7592004363e5b40ec43e1f122ed8641cd8965b
// Component : DandSocSimple
// Git hash  : 9970f6a9d3fe15fd7e1d271c3af48e12272531e8

`timescale 1ns/1ps

module DandSocSimple (
  input               io_asyncResetn,
  input               io_axiClk,
  output              io_uart_txd,
  input               io_uart_rxd
);

  wire                bufferCC_1_io_dataIn;
  wire       [31:0]   axi_downsizer_io_input_aw_payload_addr;
  wire       [3:0]    axi_downsizer_io_input_aw_payload_id;
  wire       [15:0]   axi_uartCtrl_io_apb_PADDR;
  wire                axi_uartCtrl_io_resetn;
  wire       [1:0]    core_cpu_icache_decoder_io_outputs_0_r_payload_id;
  wire       [1:0]    core_cpu_icache_decoder_io_outputs_1_r_payload_id;
  wire       [1:0]    core_cpu_dcache_decoder_io_outputs_0_r_payload_id;
  wire       [1:0]    core_cpu_dcache_decoder_io_outputs_1_r_payload_id;
  wire       [1:0]    core_cpu_dcache_decoder_1_io_outputs_0_b_payload_id;
  wire       [1:0]    core_cpu_dcache_decoder_1_io_outputs_1_b_payload_id;
  wire       [16:0]   axi_ram_io_axi_arbiter_io_readInputs_0_ar_payload_addr;
  wire       [2:0]    axi_ram_io_axi_arbiter_io_readInputs_0_ar_payload_id;
  wire       [16:0]   axi_ram_io_axi_arbiter_io_readInputs_1_ar_payload_addr;
  wire       [2:0]    axi_ram_io_axi_arbiter_io_readInputs_1_ar_payload_id;
  wire       [16:0]   axi_ram_io_axi_arbiter_io_writeInputs_0_aw_payload_addr;
  wire       [3:0]    axi_ram_io_axi_arbiter_io_writeInputs_0_aw_payload_id;
  wire       [31:0]   axi4ReadOnlyArbiter_1_io_inputs_0_ar_payload_addr;
  wire       [2:0]    axi4ReadOnlyArbiter_1_io_inputs_0_ar_payload_id;
  wire       [31:0]   axi4ReadOnlyArbiter_1_io_inputs_1_ar_payload_addr;
  wire       [2:0]    axi4ReadOnlyArbiter_1_io_inputs_1_ar_payload_id;
  wire       [16:0]   axi_bootram_io_axi_arbiter_io_readInputs_0_ar_payload_addr;
  wire       [16:0]   axi_bootram_io_axi_arbiter_io_writeInputs_0_aw_payload_addr;
  wire       [19:0]   axi_apbBridge_io_axi_arbiter_io_readInputs_0_ar_payload_addr;
  wire       [19:0]   axi_apbBridge_io_axi_arbiter_io_writeInputs_0_aw_payload_addr;
  wire                bufferCC_1_io_dataOut;
  wire                core_cpu_icache_ar_valid;
  wire       [63:0]   core_cpu_icache_ar_payload_addr;
  wire       [1:0]    core_cpu_icache_ar_payload_id;
  wire       [7:0]    core_cpu_icache_ar_payload_len;
  wire       [2:0]    core_cpu_icache_ar_payload_size;
  wire       [1:0]    core_cpu_icache_ar_payload_burst;
  wire                core_cpu_icache_r_ready;
  wire                core_cpu_dcache_ar_valid;
  wire       [63:0]   core_cpu_dcache_ar_payload_addr;
  wire       [1:0]    core_cpu_dcache_ar_payload_id;
  wire       [7:0]    core_cpu_dcache_ar_payload_len;
  wire       [2:0]    core_cpu_dcache_ar_payload_size;
  wire       [1:0]    core_cpu_dcache_ar_payload_burst;
  wire                core_cpu_dcache_r_ready;
  wire                core_cpu_dcache_aw_valid;
  wire       [63:0]   core_cpu_dcache_aw_payload_addr;
  wire       [1:0]    core_cpu_dcache_aw_payload_id;
  wire       [7:0]    core_cpu_dcache_aw_payload_len;
  wire       [2:0]    core_cpu_dcache_aw_payload_size;
  wire       [1:0]    core_cpu_dcache_aw_payload_burst;
  wire                core_cpu_dcache_w_valid;
  wire       [63:0]   core_cpu_dcache_w_payload_data;
  wire       [7:0]    core_cpu_dcache_w_payload_strb;
  wire                core_cpu_dcache_w_payload_last;
  wire                core_cpu_dcache_b_ready;
  wire                axi_downsizer_io_input_ar_ready;
  wire                axi_downsizer_io_input_aw_ready;
  wire                axi_downsizer_io_input_w_ready;
  wire                axi_downsizer_io_input_r_valid;
  wire       [63:0]   axi_downsizer_io_input_r_payload_data;
  wire       [3:0]    axi_downsizer_io_input_r_payload_id;
  wire       [1:0]    axi_downsizer_io_input_r_payload_resp;
  wire                axi_downsizer_io_input_r_payload_last;
  wire                axi_downsizer_io_input_b_valid;
  wire       [3:0]    axi_downsizer_io_input_b_payload_id;
  wire       [1:0]    axi_downsizer_io_input_b_payload_resp;
  wire                axi_downsizer_io_output_ar_valid;
  wire       [31:0]   axi_downsizer_io_output_ar_payload_addr;
  wire       [3:0]    axi_downsizer_io_output_ar_payload_id;
  wire       [3:0]    axi_downsizer_io_output_ar_payload_region;
  wire       [7:0]    axi_downsizer_io_output_ar_payload_len;
  wire       [2:0]    axi_downsizer_io_output_ar_payload_size;
  wire       [1:0]    axi_downsizer_io_output_ar_payload_burst;
  wire       [0:0]    axi_downsizer_io_output_ar_payload_lock;
  wire       [3:0]    axi_downsizer_io_output_ar_payload_cache;
  wire       [3:0]    axi_downsizer_io_output_ar_payload_qos;
  wire       [2:0]    axi_downsizer_io_output_ar_payload_prot;
  wire                axi_downsizer_io_output_aw_valid;
  wire       [31:0]   axi_downsizer_io_output_aw_payload_addr;
  wire       [3:0]    axi_downsizer_io_output_aw_payload_id;
  wire       [3:0]    axi_downsizer_io_output_aw_payload_region;
  wire       [7:0]    axi_downsizer_io_output_aw_payload_len;
  wire       [2:0]    axi_downsizer_io_output_aw_payload_size;
  wire       [1:0]    axi_downsizer_io_output_aw_payload_burst;
  wire       [0:0]    axi_downsizer_io_output_aw_payload_lock;
  wire       [3:0]    axi_downsizer_io_output_aw_payload_cache;
  wire       [3:0]    axi_downsizer_io_output_aw_payload_qos;
  wire       [2:0]    axi_downsizer_io_output_aw_payload_prot;
  wire                axi_downsizer_io_output_w_valid;
  wire       [31:0]   axi_downsizer_io_output_w_payload_data;
  wire       [3:0]    axi_downsizer_io_output_w_payload_strb;
  wire                axi_downsizer_io_output_w_payload_last;
  wire                axi_downsizer_io_output_r_ready;
  wire                axi_downsizer_io_output_b_ready;
  wire                axi_ram_io_axi_arw_ready;
  wire                axi_ram_io_axi_w_ready;
  wire                axi_ram_io_axi_b_valid;
  wire       [3:0]    axi_ram_io_axi_b_payload_id;
  wire       [1:0]    axi_ram_io_axi_b_payload_resp;
  wire                axi_ram_io_axi_r_valid;
  wire       [63:0]   axi_ram_io_axi_r_payload_data;
  wire       [3:0]    axi_ram_io_axi_r_payload_id;
  wire       [1:0]    axi_ram_io_axi_r_payload_resp;
  wire                axi_ram_io_axi_r_payload_last;
  wire                axi_bootram_io_axi_arw_ready;
  wire                axi_bootram_io_axi_w_ready;
  wire                axi_bootram_io_axi_b_valid;
  wire       [3:0]    axi_bootram_io_axi_b_payload_id;
  wire       [1:0]    axi_bootram_io_axi_b_payload_resp;
  wire                axi_bootram_io_axi_r_valid;
  wire       [31:0]   axi_bootram_io_axi_r_payload_data;
  wire       [3:0]    axi_bootram_io_axi_r_payload_id;
  wire       [1:0]    axi_bootram_io_axi_r_payload_resp;
  wire                axi_bootram_io_axi_r_payload_last;
  wire                axi_apbBridge_io_axi_arw_ready;
  wire                axi_apbBridge_io_axi_w_ready;
  wire                axi_apbBridge_io_axi_b_valid;
  wire       [3:0]    axi_apbBridge_io_axi_b_payload_id;
  wire       [1:0]    axi_apbBridge_io_axi_b_payload_resp;
  wire                axi_apbBridge_io_axi_r_valid;
  wire       [31:0]   axi_apbBridge_io_axi_r_payload_data;
  wire       [3:0]    axi_apbBridge_io_axi_r_payload_id;
  wire       [1:0]    axi_apbBridge_io_axi_r_payload_resp;
  wire                axi_apbBridge_io_axi_r_payload_last;
  wire       [19:0]   axi_apbBridge_io_apb_PADDR;
  wire       [0:0]    axi_apbBridge_io_apb_PSEL;
  wire                axi_apbBridge_io_apb_PENABLE;
  wire                axi_apbBridge_io_apb_PWRITE;
  wire       [31:0]   axi_apbBridge_io_apb_PWDATA;
  wire                axi_uartCtrl_io_apb_PREADY;
  wire       [31:0]   axi_uartCtrl_io_apb_PRDATA;
  wire                axi_uartCtrl_io_apb_PSLVERROR;
  wire                axi_uartCtrl_io_uart_txd;
  wire                core_cpu_icache_decoder_io_input_ar_ready;
  wire                core_cpu_icache_decoder_io_input_r_valid;
  wire       [63:0]   core_cpu_icache_decoder_io_input_r_payload_data;
  wire       [1:0]    core_cpu_icache_decoder_io_input_r_payload_id;
  wire       [1:0]    core_cpu_icache_decoder_io_input_r_payload_resp;
  wire                core_cpu_icache_decoder_io_input_r_payload_last;
  wire                core_cpu_icache_decoder_io_outputs_0_ar_valid;
  wire       [63:0]   core_cpu_icache_decoder_io_outputs_0_ar_payload_addr;
  wire       [1:0]    core_cpu_icache_decoder_io_outputs_0_ar_payload_id;
  wire       [7:0]    core_cpu_icache_decoder_io_outputs_0_ar_payload_len;
  wire       [2:0]    core_cpu_icache_decoder_io_outputs_0_ar_payload_size;
  wire       [1:0]    core_cpu_icache_decoder_io_outputs_0_ar_payload_burst;
  wire                core_cpu_icache_decoder_io_outputs_0_r_ready;
  wire                core_cpu_icache_decoder_io_outputs_1_ar_valid;
  wire       [63:0]   core_cpu_icache_decoder_io_outputs_1_ar_payload_addr;
  wire       [1:0]    core_cpu_icache_decoder_io_outputs_1_ar_payload_id;
  wire       [7:0]    core_cpu_icache_decoder_io_outputs_1_ar_payload_len;
  wire       [2:0]    core_cpu_icache_decoder_io_outputs_1_ar_payload_size;
  wire       [1:0]    core_cpu_icache_decoder_io_outputs_1_ar_payload_burst;
  wire                core_cpu_icache_decoder_io_outputs_1_r_ready;
  wire                core_cpu_dcache_decoder_io_input_ar_ready;
  wire                core_cpu_dcache_decoder_io_input_r_valid;
  wire       [63:0]   core_cpu_dcache_decoder_io_input_r_payload_data;
  wire       [1:0]    core_cpu_dcache_decoder_io_input_r_payload_id;
  wire       [1:0]    core_cpu_dcache_decoder_io_input_r_payload_resp;
  wire                core_cpu_dcache_decoder_io_input_r_payload_last;
  wire                core_cpu_dcache_decoder_io_outputs_0_ar_valid;
  wire       [63:0]   core_cpu_dcache_decoder_io_outputs_0_ar_payload_addr;
  wire       [1:0]    core_cpu_dcache_decoder_io_outputs_0_ar_payload_id;
  wire       [7:0]    core_cpu_dcache_decoder_io_outputs_0_ar_payload_len;
  wire       [2:0]    core_cpu_dcache_decoder_io_outputs_0_ar_payload_size;
  wire       [1:0]    core_cpu_dcache_decoder_io_outputs_0_ar_payload_burst;
  wire                core_cpu_dcache_decoder_io_outputs_0_r_ready;
  wire                core_cpu_dcache_decoder_io_outputs_1_ar_valid;
  wire       [63:0]   core_cpu_dcache_decoder_io_outputs_1_ar_payload_addr;
  wire       [1:0]    core_cpu_dcache_decoder_io_outputs_1_ar_payload_id;
  wire       [7:0]    core_cpu_dcache_decoder_io_outputs_1_ar_payload_len;
  wire       [2:0]    core_cpu_dcache_decoder_io_outputs_1_ar_payload_size;
  wire       [1:0]    core_cpu_dcache_decoder_io_outputs_1_ar_payload_burst;
  wire                core_cpu_dcache_decoder_io_outputs_1_r_ready;
  wire                core_cpu_dcache_decoder_1_io_input_aw_ready;
  wire                core_cpu_dcache_decoder_1_io_input_w_ready;
  wire                core_cpu_dcache_decoder_1_io_input_b_valid;
  wire       [1:0]    core_cpu_dcache_decoder_1_io_input_b_payload_id;
  wire       [1:0]    core_cpu_dcache_decoder_1_io_input_b_payload_resp;
  wire                core_cpu_dcache_decoder_1_io_outputs_0_aw_valid;
  wire       [63:0]   core_cpu_dcache_decoder_1_io_outputs_0_aw_payload_addr;
  wire       [1:0]    core_cpu_dcache_decoder_1_io_outputs_0_aw_payload_id;
  wire       [7:0]    core_cpu_dcache_decoder_1_io_outputs_0_aw_payload_len;
  wire       [2:0]    core_cpu_dcache_decoder_1_io_outputs_0_aw_payload_size;
  wire       [1:0]    core_cpu_dcache_decoder_1_io_outputs_0_aw_payload_burst;
  wire                core_cpu_dcache_decoder_1_io_outputs_0_w_valid;
  wire       [63:0]   core_cpu_dcache_decoder_1_io_outputs_0_w_payload_data;
  wire       [7:0]    core_cpu_dcache_decoder_1_io_outputs_0_w_payload_strb;
  wire                core_cpu_dcache_decoder_1_io_outputs_0_w_payload_last;
  wire                core_cpu_dcache_decoder_1_io_outputs_0_b_ready;
  wire                core_cpu_dcache_decoder_1_io_outputs_1_aw_valid;
  wire       [63:0]   core_cpu_dcache_decoder_1_io_outputs_1_aw_payload_addr;
  wire       [1:0]    core_cpu_dcache_decoder_1_io_outputs_1_aw_payload_id;
  wire       [7:0]    core_cpu_dcache_decoder_1_io_outputs_1_aw_payload_len;
  wire       [2:0]    core_cpu_dcache_decoder_1_io_outputs_1_aw_payload_size;
  wire       [1:0]    core_cpu_dcache_decoder_1_io_outputs_1_aw_payload_burst;
  wire                core_cpu_dcache_decoder_1_io_outputs_1_w_valid;
  wire       [63:0]   core_cpu_dcache_decoder_1_io_outputs_1_w_payload_data;
  wire       [7:0]    core_cpu_dcache_decoder_1_io_outputs_1_w_payload_strb;
  wire                core_cpu_dcache_decoder_1_io_outputs_1_w_payload_last;
  wire                core_cpu_dcache_decoder_1_io_outputs_1_b_ready;
  wire                axi_ram_io_axi_arbiter_io_readInputs_0_ar_ready;
  wire                axi_ram_io_axi_arbiter_io_readInputs_0_r_valid;
  wire       [63:0]   axi_ram_io_axi_arbiter_io_readInputs_0_r_payload_data;
  wire       [2:0]    axi_ram_io_axi_arbiter_io_readInputs_0_r_payload_id;
  wire       [1:0]    axi_ram_io_axi_arbiter_io_readInputs_0_r_payload_resp;
  wire                axi_ram_io_axi_arbiter_io_readInputs_0_r_payload_last;
  wire                axi_ram_io_axi_arbiter_io_readInputs_1_ar_ready;
  wire                axi_ram_io_axi_arbiter_io_readInputs_1_r_valid;
  wire       [63:0]   axi_ram_io_axi_arbiter_io_readInputs_1_r_payload_data;
  wire       [2:0]    axi_ram_io_axi_arbiter_io_readInputs_1_r_payload_id;
  wire       [1:0]    axi_ram_io_axi_arbiter_io_readInputs_1_r_payload_resp;
  wire                axi_ram_io_axi_arbiter_io_readInputs_1_r_payload_last;
  wire                axi_ram_io_axi_arbiter_io_writeInputs_0_aw_ready;
  wire                axi_ram_io_axi_arbiter_io_writeInputs_0_w_ready;
  wire                axi_ram_io_axi_arbiter_io_writeInputs_0_b_valid;
  wire       [3:0]    axi_ram_io_axi_arbiter_io_writeInputs_0_b_payload_id;
  wire       [1:0]    axi_ram_io_axi_arbiter_io_writeInputs_0_b_payload_resp;
  wire                axi_ram_io_axi_arbiter_io_output_arw_valid;
  wire       [16:0]   axi_ram_io_axi_arbiter_io_output_arw_payload_addr;
  wire       [3:0]    axi_ram_io_axi_arbiter_io_output_arw_payload_id;
  wire       [7:0]    axi_ram_io_axi_arbiter_io_output_arw_payload_len;
  wire       [2:0]    axi_ram_io_axi_arbiter_io_output_arw_payload_size;
  wire       [1:0]    axi_ram_io_axi_arbiter_io_output_arw_payload_burst;
  wire                axi_ram_io_axi_arbiter_io_output_arw_payload_write;
  wire                axi_ram_io_axi_arbiter_io_output_w_valid;
  wire       [63:0]   axi_ram_io_axi_arbiter_io_output_w_payload_data;
  wire       [7:0]    axi_ram_io_axi_arbiter_io_output_w_payload_strb;
  wire                axi_ram_io_axi_arbiter_io_output_w_payload_last;
  wire                axi_ram_io_axi_arbiter_io_output_b_ready;
  wire                axi_ram_io_axi_arbiter_io_output_r_ready;
  wire                axi4ReadOnlyArbiter_1_io_inputs_0_ar_ready;
  wire                axi4ReadOnlyArbiter_1_io_inputs_0_r_valid;
  wire       [63:0]   axi4ReadOnlyArbiter_1_io_inputs_0_r_payload_data;
  wire       [2:0]    axi4ReadOnlyArbiter_1_io_inputs_0_r_payload_id;
  wire       [1:0]    axi4ReadOnlyArbiter_1_io_inputs_0_r_payload_resp;
  wire                axi4ReadOnlyArbiter_1_io_inputs_0_r_payload_last;
  wire                axi4ReadOnlyArbiter_1_io_inputs_1_ar_ready;
  wire                axi4ReadOnlyArbiter_1_io_inputs_1_r_valid;
  wire       [63:0]   axi4ReadOnlyArbiter_1_io_inputs_1_r_payload_data;
  wire       [2:0]    axi4ReadOnlyArbiter_1_io_inputs_1_r_payload_id;
  wire       [1:0]    axi4ReadOnlyArbiter_1_io_inputs_1_r_payload_resp;
  wire                axi4ReadOnlyArbiter_1_io_inputs_1_r_payload_last;
  wire                axi4ReadOnlyArbiter_1_io_output_ar_valid;
  wire       [31:0]   axi4ReadOnlyArbiter_1_io_output_ar_payload_addr;
  wire       [3:0]    axi4ReadOnlyArbiter_1_io_output_ar_payload_id;
  wire       [3:0]    axi4ReadOnlyArbiter_1_io_output_ar_payload_region;
  wire       [7:0]    axi4ReadOnlyArbiter_1_io_output_ar_payload_len;
  wire       [2:0]    axi4ReadOnlyArbiter_1_io_output_ar_payload_size;
  wire       [1:0]    axi4ReadOnlyArbiter_1_io_output_ar_payload_burst;
  wire       [0:0]    axi4ReadOnlyArbiter_1_io_output_ar_payload_lock;
  wire       [3:0]    axi4ReadOnlyArbiter_1_io_output_ar_payload_cache;
  wire       [3:0]    axi4ReadOnlyArbiter_1_io_output_ar_payload_qos;
  wire       [2:0]    axi4ReadOnlyArbiter_1_io_output_ar_payload_prot;
  wire                axi4ReadOnlyArbiter_1_io_output_r_ready;
  wire                toplevel_axi_downsizer_io_output_readOnly_decoder_io_input_ar_ready;
  wire                toplevel_axi_downsizer_io_output_readOnly_decoder_io_input_r_valid;
  wire       [31:0]   toplevel_axi_downsizer_io_output_readOnly_decoder_io_input_r_payload_data;
  wire       [3:0]    toplevel_axi_downsizer_io_output_readOnly_decoder_io_input_r_payload_id;
  wire       [1:0]    toplevel_axi_downsizer_io_output_readOnly_decoder_io_input_r_payload_resp;
  wire                toplevel_axi_downsizer_io_output_readOnly_decoder_io_input_r_payload_last;
  wire                toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_valid;
  wire       [31:0]   toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_payload_addr;
  wire       [3:0]    toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_payload_id;
  wire       [3:0]    toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_payload_region;
  wire       [7:0]    toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_payload_len;
  wire       [2:0]    toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_payload_size;
  wire       [1:0]    toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_payload_burst;
  wire       [0:0]    toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_payload_lock;
  wire       [3:0]    toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_payload_cache;
  wire       [3:0]    toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_payload_qos;
  wire       [2:0]    toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_payload_prot;
  wire                toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_r_ready;
  wire                toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_valid;
  wire       [31:0]   toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_payload_addr;
  wire       [3:0]    toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_payload_id;
  wire       [3:0]    toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_payload_region;
  wire       [7:0]    toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_payload_len;
  wire       [2:0]    toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_payload_size;
  wire       [1:0]    toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_payload_burst;
  wire       [0:0]    toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_payload_lock;
  wire       [3:0]    toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_payload_cache;
  wire       [3:0]    toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_payload_qos;
  wire       [2:0]    toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_payload_prot;
  wire                toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_r_ready;
  wire                toplevel_axi_downsizer_io_output_writeOnly_decoder_io_input_aw_ready;
  wire                toplevel_axi_downsizer_io_output_writeOnly_decoder_io_input_w_ready;
  wire                toplevel_axi_downsizer_io_output_writeOnly_decoder_io_input_b_valid;
  wire       [3:0]    toplevel_axi_downsizer_io_output_writeOnly_decoder_io_input_b_payload_id;
  wire       [1:0]    toplevel_axi_downsizer_io_output_writeOnly_decoder_io_input_b_payload_resp;
  wire                toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_valid;
  wire       [31:0]   toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_payload_addr;
  wire       [3:0]    toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_payload_id;
  wire       [3:0]    toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_payload_region;
  wire       [7:0]    toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_payload_len;
  wire       [2:0]    toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_payload_size;
  wire       [1:0]    toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_payload_burst;
  wire       [0:0]    toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_payload_lock;
  wire       [3:0]    toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_payload_cache;
  wire       [3:0]    toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_payload_qos;
  wire       [2:0]    toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_payload_prot;
  wire                toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_w_valid;
  wire       [31:0]   toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_w_payload_data;
  wire       [3:0]    toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_w_payload_strb;
  wire                toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_w_payload_last;
  wire                toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_b_ready;
  wire                toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_valid;
  wire       [31:0]   toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_payload_addr;
  wire       [3:0]    toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_payload_id;
  wire       [3:0]    toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_payload_region;
  wire       [7:0]    toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_payload_len;
  wire       [2:0]    toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_payload_size;
  wire       [1:0]    toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_payload_burst;
  wire       [0:0]    toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_payload_lock;
  wire       [3:0]    toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_payload_cache;
  wire       [3:0]    toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_payload_qos;
  wire       [2:0]    toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_payload_prot;
  wire                toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_w_valid;
  wire       [31:0]   toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_w_payload_data;
  wire       [3:0]    toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_w_payload_strb;
  wire                toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_w_payload_last;
  wire                toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_b_ready;
  wire                axi_bootram_io_axi_arbiter_io_readInputs_0_ar_ready;
  wire                axi_bootram_io_axi_arbiter_io_readInputs_0_r_valid;
  wire       [31:0]   axi_bootram_io_axi_arbiter_io_readInputs_0_r_payload_data;
  wire       [3:0]    axi_bootram_io_axi_arbiter_io_readInputs_0_r_payload_id;
  wire       [1:0]    axi_bootram_io_axi_arbiter_io_readInputs_0_r_payload_resp;
  wire                axi_bootram_io_axi_arbiter_io_readInputs_0_r_payload_last;
  wire                axi_bootram_io_axi_arbiter_io_writeInputs_0_aw_ready;
  wire                axi_bootram_io_axi_arbiter_io_writeInputs_0_w_ready;
  wire                axi_bootram_io_axi_arbiter_io_writeInputs_0_b_valid;
  wire       [3:0]    axi_bootram_io_axi_arbiter_io_writeInputs_0_b_payload_id;
  wire       [1:0]    axi_bootram_io_axi_arbiter_io_writeInputs_0_b_payload_resp;
  wire                axi_bootram_io_axi_arbiter_io_output_arw_valid;
  wire       [16:0]   axi_bootram_io_axi_arbiter_io_output_arw_payload_addr;
  wire       [3:0]    axi_bootram_io_axi_arbiter_io_output_arw_payload_id;
  wire       [7:0]    axi_bootram_io_axi_arbiter_io_output_arw_payload_len;
  wire       [2:0]    axi_bootram_io_axi_arbiter_io_output_arw_payload_size;
  wire       [1:0]    axi_bootram_io_axi_arbiter_io_output_arw_payload_burst;
  wire                axi_bootram_io_axi_arbiter_io_output_arw_payload_write;
  wire                axi_bootram_io_axi_arbiter_io_output_w_valid;
  wire       [31:0]   axi_bootram_io_axi_arbiter_io_output_w_payload_data;
  wire       [3:0]    axi_bootram_io_axi_arbiter_io_output_w_payload_strb;
  wire                axi_bootram_io_axi_arbiter_io_output_w_payload_last;
  wire                axi_bootram_io_axi_arbiter_io_output_b_ready;
  wire                axi_bootram_io_axi_arbiter_io_output_r_ready;
  wire                axi_apbBridge_io_axi_arbiter_io_readInputs_0_ar_ready;
  wire                axi_apbBridge_io_axi_arbiter_io_readInputs_0_r_valid;
  wire       [31:0]   axi_apbBridge_io_axi_arbiter_io_readInputs_0_r_payload_data;
  wire       [3:0]    axi_apbBridge_io_axi_arbiter_io_readInputs_0_r_payload_id;
  wire       [1:0]    axi_apbBridge_io_axi_arbiter_io_readInputs_0_r_payload_resp;
  wire                axi_apbBridge_io_axi_arbiter_io_readInputs_0_r_payload_last;
  wire                axi_apbBridge_io_axi_arbiter_io_writeInputs_0_aw_ready;
  wire                axi_apbBridge_io_axi_arbiter_io_writeInputs_0_w_ready;
  wire                axi_apbBridge_io_axi_arbiter_io_writeInputs_0_b_valid;
  wire       [3:0]    axi_apbBridge_io_axi_arbiter_io_writeInputs_0_b_payload_id;
  wire       [1:0]    axi_apbBridge_io_axi_arbiter_io_writeInputs_0_b_payload_resp;
  wire                axi_apbBridge_io_axi_arbiter_io_output_arw_valid;
  wire       [19:0]   axi_apbBridge_io_axi_arbiter_io_output_arw_payload_addr;
  wire       [3:0]    axi_apbBridge_io_axi_arbiter_io_output_arw_payload_id;
  wire       [7:0]    axi_apbBridge_io_axi_arbiter_io_output_arw_payload_len;
  wire       [2:0]    axi_apbBridge_io_axi_arbiter_io_output_arw_payload_size;
  wire       [1:0]    axi_apbBridge_io_axi_arbiter_io_output_arw_payload_burst;
  wire                axi_apbBridge_io_axi_arbiter_io_output_arw_payload_write;
  wire                axi_apbBridge_io_axi_arbiter_io_output_w_valid;
  wire       [31:0]   axi_apbBridge_io_axi_arbiter_io_output_w_payload_data;
  wire       [3:0]    axi_apbBridge_io_axi_arbiter_io_output_w_payload_strb;
  wire                axi_apbBridge_io_axi_arbiter_io_output_w_payload_last;
  wire                axi_apbBridge_io_axi_arbiter_io_output_b_ready;
  wire                axi_apbBridge_io_axi_arbiter_io_output_r_ready;
  wire                io_apb_decoder_io_input_PREADY;
  wire       [31:0]   io_apb_decoder_io_input_PRDATA;
  wire                io_apb_decoder_io_input_PSLVERROR;
  wire       [19:0]   io_apb_decoder_io_output_PADDR;
  wire       [0:0]    io_apb_decoder_io_output_PSEL;
  wire                io_apb_decoder_io_output_PENABLE;
  wire                io_apb_decoder_io_output_PWRITE;
  wire       [31:0]   io_apb_decoder_io_output_PWDATA;
  wire                apb3Router_1_io_input_PREADY;
  wire       [31:0]   apb3Router_1_io_input_PRDATA;
  wire                apb3Router_1_io_input_PSLVERROR;
  wire       [19:0]   apb3Router_1_io_outputs_0_PADDR;
  wire       [0:0]    apb3Router_1_io_outputs_0_PSEL;
  wire                apb3Router_1_io_outputs_0_PENABLE;
  wire                apb3Router_1_io_outputs_0_PWRITE;
  wire       [31:0]   apb3Router_1_io_outputs_0_PWDATA;
  reg                 resetCtrl_systemResetUnbuffered;
  reg        [5:0]    resetCtrl_systemResetCounter;
  wire       [5:0]    _zz_when_GenDandSocSimple_l89;
  wire                when_GenDandSocSimple_l89;
  wire                when_GenDandSocSimple_l93;
  reg                 resetCtrl_axiReset;
  wire                toplevel_axi_downsizer_io_output_readOnly_ar_valid;
  wire                toplevel_axi_downsizer_io_output_readOnly_ar_ready;
  wire       [31:0]   toplevel_axi_downsizer_io_output_readOnly_ar_payload_addr;
  wire       [3:0]    toplevel_axi_downsizer_io_output_readOnly_ar_payload_id;
  wire       [3:0]    toplevel_axi_downsizer_io_output_readOnly_ar_payload_region;
  wire       [7:0]    toplevel_axi_downsizer_io_output_readOnly_ar_payload_len;
  wire       [2:0]    toplevel_axi_downsizer_io_output_readOnly_ar_payload_size;
  wire       [1:0]    toplevel_axi_downsizer_io_output_readOnly_ar_payload_burst;
  wire       [0:0]    toplevel_axi_downsizer_io_output_readOnly_ar_payload_lock;
  wire       [3:0]    toplevel_axi_downsizer_io_output_readOnly_ar_payload_cache;
  wire       [3:0]    toplevel_axi_downsizer_io_output_readOnly_ar_payload_qos;
  wire       [2:0]    toplevel_axi_downsizer_io_output_readOnly_ar_payload_prot;
  wire                toplevel_axi_downsizer_io_output_readOnly_r_valid;
  wire                toplevel_axi_downsizer_io_output_readOnly_r_ready;
  wire       [31:0]   toplevel_axi_downsizer_io_output_readOnly_r_payload_data;
  wire       [3:0]    toplevel_axi_downsizer_io_output_readOnly_r_payload_id;
  wire       [1:0]    toplevel_axi_downsizer_io_output_readOnly_r_payload_resp;
  wire                toplevel_axi_downsizer_io_output_readOnly_r_payload_last;
  wire                toplevel_axi_downsizer_io_output_writeOnly_aw_valid;
  wire                toplevel_axi_downsizer_io_output_writeOnly_aw_ready;
  wire       [31:0]   toplevel_axi_downsizer_io_output_writeOnly_aw_payload_addr;
  wire       [3:0]    toplevel_axi_downsizer_io_output_writeOnly_aw_payload_id;
  wire       [3:0]    toplevel_axi_downsizer_io_output_writeOnly_aw_payload_region;
  wire       [7:0]    toplevel_axi_downsizer_io_output_writeOnly_aw_payload_len;
  wire       [2:0]    toplevel_axi_downsizer_io_output_writeOnly_aw_payload_size;
  wire       [1:0]    toplevel_axi_downsizer_io_output_writeOnly_aw_payload_burst;
  wire       [0:0]    toplevel_axi_downsizer_io_output_writeOnly_aw_payload_lock;
  wire       [3:0]    toplevel_axi_downsizer_io_output_writeOnly_aw_payload_cache;
  wire       [3:0]    toplevel_axi_downsizer_io_output_writeOnly_aw_payload_qos;
  wire       [2:0]    toplevel_axi_downsizer_io_output_writeOnly_aw_payload_prot;
  wire                toplevel_axi_downsizer_io_output_writeOnly_w_valid;
  wire                toplevel_axi_downsizer_io_output_writeOnly_w_ready;
  wire       [31:0]   toplevel_axi_downsizer_io_output_writeOnly_w_payload_data;
  wire       [3:0]    toplevel_axi_downsizer_io_output_writeOnly_w_payload_strb;
  wire                toplevel_axi_downsizer_io_output_writeOnly_w_payload_last;
  wire                toplevel_axi_downsizer_io_output_writeOnly_b_valid;
  wire                toplevel_axi_downsizer_io_output_writeOnly_b_ready;
  wire       [3:0]    toplevel_axi_downsizer_io_output_writeOnly_b_payload_id;
  wire       [1:0]    toplevel_axi_downsizer_io_output_writeOnly_b_payload_resp;
  wire                toplevel_core_cpu_icache_decoder_io_outputs_0_ar_validPipe_valid;
  wire                toplevel_core_cpu_icache_decoder_io_outputs_0_ar_validPipe_ready;
  wire       [63:0]   toplevel_core_cpu_icache_decoder_io_outputs_0_ar_validPipe_payload_addr;
  wire       [1:0]    toplevel_core_cpu_icache_decoder_io_outputs_0_ar_validPipe_payload_id;
  wire       [7:0]    toplevel_core_cpu_icache_decoder_io_outputs_0_ar_validPipe_payload_len;
  wire       [2:0]    toplevel_core_cpu_icache_decoder_io_outputs_0_ar_validPipe_payload_size;
  wire       [1:0]    toplevel_core_cpu_icache_decoder_io_outputs_0_ar_validPipe_payload_burst;
  reg                 toplevel_core_cpu_icache_decoder_io_outputs_0_ar_rValid;
  wire                toplevel_core_cpu_icache_decoder_io_outputs_0_ar_validPipe_fire;
  wire                toplevel_core_cpu_icache_decoder_io_outputs_0_ar_validPipe_fire_1;
  wire                toplevel_core_cpu_icache_decoder_io_outputs_1_ar_validPipe_valid;
  wire                toplevel_core_cpu_icache_decoder_io_outputs_1_ar_validPipe_ready;
  wire       [63:0]   toplevel_core_cpu_icache_decoder_io_outputs_1_ar_validPipe_payload_addr;
  wire       [1:0]    toplevel_core_cpu_icache_decoder_io_outputs_1_ar_validPipe_payload_id;
  wire       [7:0]    toplevel_core_cpu_icache_decoder_io_outputs_1_ar_validPipe_payload_len;
  wire       [2:0]    toplevel_core_cpu_icache_decoder_io_outputs_1_ar_validPipe_payload_size;
  wire       [1:0]    toplevel_core_cpu_icache_decoder_io_outputs_1_ar_validPipe_payload_burst;
  reg                 toplevel_core_cpu_icache_decoder_io_outputs_1_ar_rValid;
  wire                toplevel_core_cpu_icache_decoder_io_outputs_1_ar_validPipe_fire;
  wire                toplevel_core_cpu_icache_decoder_io_outputs_1_ar_validPipe_fire_1;
  wire                toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_validPipe_valid;
  wire                toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_validPipe_ready;
  wire       [63:0]   toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_validPipe_payload_addr;
  wire       [1:0]    toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_validPipe_payload_id;
  wire       [7:0]    toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_validPipe_payload_len;
  wire       [2:0]    toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_validPipe_payload_size;
  wire       [1:0]    toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_validPipe_payload_burst;
  reg                 toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_rValid;
  wire                toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_validPipe_fire;
  wire                toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_validPipe_fire_1;
  wire                toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_validPipe_valid;
  wire                toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_validPipe_ready;
  wire       [63:0]   toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_validPipe_payload_addr;
  wire       [1:0]    toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_validPipe_payload_id;
  wire       [7:0]    toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_validPipe_payload_len;
  wire       [2:0]    toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_validPipe_payload_size;
  wire       [1:0]    toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_validPipe_payload_burst;
  reg                 toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_rValid;
  wire                toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_validPipe_fire;
  wire                toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_validPipe_fire_1;
  wire                toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_validPipe_valid;
  wire                toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_validPipe_ready;
  wire       [63:0]   toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_validPipe_payload_addr;
  wire       [1:0]    toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_validPipe_payload_id;
  wire       [7:0]    toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_validPipe_payload_len;
  wire       [2:0]    toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_validPipe_payload_size;
  wire       [1:0]    toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_validPipe_payload_burst;
  reg                 toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_rValid;
  wire                toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_validPipe_fire;
  wire                toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_validPipe_fire_1;
  wire                toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_validPipe_valid;
  wire                toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_validPipe_ready;
  wire       [63:0]   toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_validPipe_payload_addr;
  wire       [1:0]    toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_validPipe_payload_id;
  wire       [7:0]    toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_validPipe_payload_len;
  wire       [2:0]    toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_validPipe_payload_size;
  wire       [1:0]    toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_validPipe_payload_burst;
  reg                 toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_rValid;
  wire                toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_validPipe_fire;
  wire                toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_validPipe_fire_1;
  wire       [3:0]    _zz_io_inputs_0_ar_payload_region;
  wire       [3:0]    _zz_io_inputs_1_ar_payload_region;
  wire       [3:0]    _zz_io_input_aw_payload_region;
  wire                toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_valid;
  wire                toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_ready;
  wire       [31:0]   toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_payload_addr;
  wire       [3:0]    toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_payload_id;
  wire       [3:0]    toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_payload_region;
  wire       [7:0]    toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_payload_len;
  wire       [2:0]    toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_payload_size;
  wire       [1:0]    toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_payload_burst;
  wire       [0:0]    toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_payload_lock;
  wire       [3:0]    toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_payload_cache;
  wire       [3:0]    toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_payload_qos;
  wire       [2:0]    toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_payload_prot;
  reg                 toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_rValid;
  wire                toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_fire;
  wire                toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_fire_1;
  wire                toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_valid;
  wire                toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_ready;
  wire       [31:0]   toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_payload_addr;
  wire       [3:0]    toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_payload_id;
  wire       [3:0]    toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_payload_region;
  wire       [7:0]    toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_payload_len;
  wire       [2:0]    toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_payload_size;
  wire       [1:0]    toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_payload_burst;
  wire       [0:0]    toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_payload_lock;
  wire       [3:0]    toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_payload_cache;
  wire       [3:0]    toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_payload_qos;
  wire       [2:0]    toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_payload_prot;
  reg                 toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_rValid;
  wire                toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_fire;
  wire                toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_fire_1;
  wire                toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_valid;
  wire                toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_ready;
  wire       [31:0]   toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_addr;
  wire       [3:0]    toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_id;
  wire       [3:0]    toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_region;
  wire       [7:0]    toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_len;
  wire       [2:0]    toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_size;
  wire       [1:0]    toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_burst;
  wire       [0:0]    toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_lock;
  wire       [3:0]    toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_cache;
  wire       [3:0]    toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_qos;
  wire       [2:0]    toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_prot;
  reg                 toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_rValid;
  wire                toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_fire;
  wire                toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_fire_1;
  wire                toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_valid;
  wire                toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_ready;
  wire       [31:0]   toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_payload_addr;
  wire       [3:0]    toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_payload_id;
  wire       [3:0]    toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_payload_region;
  wire       [7:0]    toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_payload_len;
  wire       [2:0]    toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_payload_size;
  wire       [1:0]    toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_payload_burst;
  wire       [0:0]    toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_payload_lock;
  wire       [3:0]    toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_payload_cache;
  wire       [3:0]    toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_payload_qos;
  wire       [2:0]    toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_payload_prot;
  reg                 toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_rValid;
  wire                toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_fire;
  wire                toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_fire_1;

  BufferCC bufferCC_1 (
    .io_dataIn      (bufferCC_1_io_dataIn ), //i
    .io_dataOut     (bufferCC_1_io_dataOut), //o
    .io_axiClk      (io_axiClk            ), //i
    .io_asyncResetn (io_asyncResetn       )  //i
  );
  DandRiscvSimple core_cpu (
    .icache_ar_valid         (core_cpu_icache_ar_valid                              ), //o
    .icache_ar_ready         (core_cpu_icache_decoder_io_input_ar_ready             ), //i
    .icache_ar_payload_addr  (core_cpu_icache_ar_payload_addr[63:0]                 ), //o
    .icache_ar_payload_id    (core_cpu_icache_ar_payload_id[1:0]                    ), //o
    .icache_ar_payload_len   (core_cpu_icache_ar_payload_len[7:0]                   ), //o
    .icache_ar_payload_size  (core_cpu_icache_ar_payload_size[2:0]                  ), //o
    .icache_ar_payload_burst (core_cpu_icache_ar_payload_burst[1:0]                 ), //o
    .icache_r_valid          (core_cpu_icache_decoder_io_input_r_valid              ), //i
    .icache_r_ready          (core_cpu_icache_r_ready                               ), //o
    .icache_r_payload_data   (core_cpu_icache_decoder_io_input_r_payload_data[63:0] ), //i
    .icache_r_payload_id     (core_cpu_icache_decoder_io_input_r_payload_id[1:0]    ), //i
    .icache_r_payload_resp   (core_cpu_icache_decoder_io_input_r_payload_resp[1:0]  ), //i
    .icache_r_payload_last   (core_cpu_icache_decoder_io_input_r_payload_last       ), //i
    .dcache_ar_valid         (core_cpu_dcache_ar_valid                              ), //o
    .dcache_ar_ready         (core_cpu_dcache_decoder_io_input_ar_ready             ), //i
    .dcache_ar_payload_addr  (core_cpu_dcache_ar_payload_addr[63:0]                 ), //o
    .dcache_ar_payload_id    (core_cpu_dcache_ar_payload_id[1:0]                    ), //o
    .dcache_ar_payload_len   (core_cpu_dcache_ar_payload_len[7:0]                   ), //o
    .dcache_ar_payload_size  (core_cpu_dcache_ar_payload_size[2:0]                  ), //o
    .dcache_ar_payload_burst (core_cpu_dcache_ar_payload_burst[1:0]                 ), //o
    .dcache_r_valid          (core_cpu_dcache_decoder_io_input_r_valid              ), //i
    .dcache_r_ready          (core_cpu_dcache_r_ready                               ), //o
    .dcache_r_payload_data   (core_cpu_dcache_decoder_io_input_r_payload_data[63:0] ), //i
    .dcache_r_payload_id     (core_cpu_dcache_decoder_io_input_r_payload_id[1:0]    ), //i
    .dcache_r_payload_resp   (core_cpu_dcache_decoder_io_input_r_payload_resp[1:0]  ), //i
    .dcache_r_payload_last   (core_cpu_dcache_decoder_io_input_r_payload_last       ), //i
    .dcache_aw_valid         (core_cpu_dcache_aw_valid                              ), //o
    .dcache_aw_ready         (core_cpu_dcache_decoder_1_io_input_aw_ready           ), //i
    .dcache_aw_payload_addr  (core_cpu_dcache_aw_payload_addr[63:0]                 ), //o
    .dcache_aw_payload_id    (core_cpu_dcache_aw_payload_id[1:0]                    ), //o
    .dcache_aw_payload_len   (core_cpu_dcache_aw_payload_len[7:0]                   ), //o
    .dcache_aw_payload_size  (core_cpu_dcache_aw_payload_size[2:0]                  ), //o
    .dcache_aw_payload_burst (core_cpu_dcache_aw_payload_burst[1:0]                 ), //o
    .dcache_w_valid          (core_cpu_dcache_w_valid                               ), //o
    .dcache_w_ready          (core_cpu_dcache_decoder_1_io_input_w_ready            ), //i
    .dcache_w_payload_data   (core_cpu_dcache_w_payload_data[63:0]                  ), //o
    .dcache_w_payload_strb   (core_cpu_dcache_w_payload_strb[7:0]                   ), //o
    .dcache_w_payload_last   (core_cpu_dcache_w_payload_last                        ), //o
    .dcache_b_valid          (core_cpu_dcache_decoder_1_io_input_b_valid            ), //i
    .dcache_b_ready          (core_cpu_dcache_b_ready                               ), //o
    .dcache_b_payload_id     (core_cpu_dcache_decoder_1_io_input_b_payload_id[1:0]  ), //i
    .dcache_b_payload_resp   (core_cpu_dcache_decoder_1_io_input_b_payload_resp[1:0]), //i
    .io_axiClk               (io_axiClk                                             ), //i
    .resetCtrl_axiReset      (resetCtrl_axiReset                                    )  //i
  );
  Axi4Downsizer axi_downsizer (
    .io_input_aw_valid           (toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_validPipe_valid             ), //i
    .io_input_aw_ready           (axi_downsizer_io_input_aw_ready                                                ), //o
    .io_input_aw_payload_addr    (axi_downsizer_io_input_aw_payload_addr[31:0]                                   ), //i
    .io_input_aw_payload_id      (axi_downsizer_io_input_aw_payload_id[3:0]                                      ), //i
    .io_input_aw_payload_region  (_zz_io_input_aw_payload_region[3:0]                                            ), //i
    .io_input_aw_payload_len     (toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_validPipe_payload_len[7:0]  ), //i
    .io_input_aw_payload_size    (toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_validPipe_payload_size[2:0] ), //i
    .io_input_aw_payload_burst   (toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_validPipe_payload_burst[1:0]), //i
    .io_input_aw_payload_lock    (1'b0                                                                           ), //i
    .io_input_aw_payload_cache   (4'b0000                                                                        ), //i
    .io_input_aw_payload_qos     (4'b0000                                                                        ), //i
    .io_input_aw_payload_prot    (3'b010                                                                         ), //i
    .io_input_w_valid            (core_cpu_dcache_decoder_1_io_outputs_1_w_valid                                 ), //i
    .io_input_w_ready            (axi_downsizer_io_input_w_ready                                                 ), //o
    .io_input_w_payload_data     (core_cpu_dcache_decoder_1_io_outputs_1_w_payload_data[63:0]                    ), //i
    .io_input_w_payload_strb     (core_cpu_dcache_decoder_1_io_outputs_1_w_payload_strb[7:0]                     ), //i
    .io_input_w_payload_last     (core_cpu_dcache_decoder_1_io_outputs_1_w_payload_last                          ), //i
    .io_input_b_valid            (axi_downsizer_io_input_b_valid                                                 ), //o
    .io_input_b_ready            (core_cpu_dcache_decoder_1_io_outputs_1_b_ready                                 ), //i
    .io_input_b_payload_id       (axi_downsizer_io_input_b_payload_id[3:0]                                       ), //o
    .io_input_b_payload_resp     (axi_downsizer_io_input_b_payload_resp[1:0]                                     ), //o
    .io_input_ar_valid           (axi4ReadOnlyArbiter_1_io_output_ar_valid                                       ), //i
    .io_input_ar_ready           (axi_downsizer_io_input_ar_ready                                                ), //o
    .io_input_ar_payload_addr    (axi4ReadOnlyArbiter_1_io_output_ar_payload_addr[31:0]                          ), //i
    .io_input_ar_payload_id      (axi4ReadOnlyArbiter_1_io_output_ar_payload_id[3:0]                             ), //i
    .io_input_ar_payload_region  (axi4ReadOnlyArbiter_1_io_output_ar_payload_region[3:0]                         ), //i
    .io_input_ar_payload_len     (axi4ReadOnlyArbiter_1_io_output_ar_payload_len[7:0]                            ), //i
    .io_input_ar_payload_size    (axi4ReadOnlyArbiter_1_io_output_ar_payload_size[2:0]                           ), //i
    .io_input_ar_payload_burst   (axi4ReadOnlyArbiter_1_io_output_ar_payload_burst[1:0]                          ), //i
    .io_input_ar_payload_lock    (axi4ReadOnlyArbiter_1_io_output_ar_payload_lock                                ), //i
    .io_input_ar_payload_cache   (axi4ReadOnlyArbiter_1_io_output_ar_payload_cache[3:0]                          ), //i
    .io_input_ar_payload_qos     (axi4ReadOnlyArbiter_1_io_output_ar_payload_qos[3:0]                            ), //i
    .io_input_ar_payload_prot    (axi4ReadOnlyArbiter_1_io_output_ar_payload_prot[2:0]                           ), //i
    .io_input_r_valid            (axi_downsizer_io_input_r_valid                                                 ), //o
    .io_input_r_ready            (axi4ReadOnlyArbiter_1_io_output_r_ready                                        ), //i
    .io_input_r_payload_data     (axi_downsizer_io_input_r_payload_data[63:0]                                    ), //o
    .io_input_r_payload_id       (axi_downsizer_io_input_r_payload_id[3:0]                                       ), //o
    .io_input_r_payload_resp     (axi_downsizer_io_input_r_payload_resp[1:0]                                     ), //o
    .io_input_r_payload_last     (axi_downsizer_io_input_r_payload_last                                          ), //o
    .io_output_aw_valid          (axi_downsizer_io_output_aw_valid                                               ), //o
    .io_output_aw_ready          (toplevel_axi_downsizer_io_output_writeOnly_aw_ready                            ), //i
    .io_output_aw_payload_addr   (axi_downsizer_io_output_aw_payload_addr[31:0]                                  ), //o
    .io_output_aw_payload_id     (axi_downsizer_io_output_aw_payload_id[3:0]                                     ), //o
    .io_output_aw_payload_region (axi_downsizer_io_output_aw_payload_region[3:0]                                 ), //o
    .io_output_aw_payload_len    (axi_downsizer_io_output_aw_payload_len[7:0]                                    ), //o
    .io_output_aw_payload_size   (axi_downsizer_io_output_aw_payload_size[2:0]                                   ), //o
    .io_output_aw_payload_burst  (axi_downsizer_io_output_aw_payload_burst[1:0]                                  ), //o
    .io_output_aw_payload_lock   (axi_downsizer_io_output_aw_payload_lock                                        ), //o
    .io_output_aw_payload_cache  (axi_downsizer_io_output_aw_payload_cache[3:0]                                  ), //o
    .io_output_aw_payload_qos    (axi_downsizer_io_output_aw_payload_qos[3:0]                                    ), //o
    .io_output_aw_payload_prot   (axi_downsizer_io_output_aw_payload_prot[2:0]                                   ), //o
    .io_output_w_valid           (axi_downsizer_io_output_w_valid                                                ), //o
    .io_output_w_ready           (toplevel_axi_downsizer_io_output_writeOnly_w_ready                             ), //i
    .io_output_w_payload_data    (axi_downsizer_io_output_w_payload_data[31:0]                                   ), //o
    .io_output_w_payload_strb    (axi_downsizer_io_output_w_payload_strb[3:0]                                    ), //o
    .io_output_w_payload_last    (axi_downsizer_io_output_w_payload_last                                         ), //o
    .io_output_b_valid           (toplevel_axi_downsizer_io_output_writeOnly_b_valid                             ), //i
    .io_output_b_ready           (axi_downsizer_io_output_b_ready                                                ), //o
    .io_output_b_payload_id      (toplevel_axi_downsizer_io_output_writeOnly_b_payload_id[3:0]                   ), //i
    .io_output_b_payload_resp    (toplevel_axi_downsizer_io_output_writeOnly_b_payload_resp[1:0]                 ), //i
    .io_output_ar_valid          (axi_downsizer_io_output_ar_valid                                               ), //o
    .io_output_ar_ready          (toplevel_axi_downsizer_io_output_readOnly_ar_ready                             ), //i
    .io_output_ar_payload_addr   (axi_downsizer_io_output_ar_payload_addr[31:0]                                  ), //o
    .io_output_ar_payload_id     (axi_downsizer_io_output_ar_payload_id[3:0]                                     ), //o
    .io_output_ar_payload_region (axi_downsizer_io_output_ar_payload_region[3:0]                                 ), //o
    .io_output_ar_payload_len    (axi_downsizer_io_output_ar_payload_len[7:0]                                    ), //o
    .io_output_ar_payload_size   (axi_downsizer_io_output_ar_payload_size[2:0]                                   ), //o
    .io_output_ar_payload_burst  (axi_downsizer_io_output_ar_payload_burst[1:0]                                  ), //o
    .io_output_ar_payload_lock   (axi_downsizer_io_output_ar_payload_lock                                        ), //o
    .io_output_ar_payload_cache  (axi_downsizer_io_output_ar_payload_cache[3:0]                                  ), //o
    .io_output_ar_payload_qos    (axi_downsizer_io_output_ar_payload_qos[3:0]                                    ), //o
    .io_output_ar_payload_prot   (axi_downsizer_io_output_ar_payload_prot[2:0]                                   ), //o
    .io_output_r_valid           (toplevel_axi_downsizer_io_output_readOnly_r_valid                              ), //i
    .io_output_r_ready           (axi_downsizer_io_output_r_ready                                                ), //o
    .io_output_r_payload_data    (toplevel_axi_downsizer_io_output_readOnly_r_payload_data[31:0]                 ), //i
    .io_output_r_payload_id      (toplevel_axi_downsizer_io_output_readOnly_r_payload_id[3:0]                    ), //i
    .io_output_r_payload_resp    (toplevel_axi_downsizer_io_output_readOnly_r_payload_resp[1:0]                  ), //i
    .io_output_r_payload_last    (toplevel_axi_downsizer_io_output_readOnly_r_payload_last                       ), //i
    .io_axiClk                   (io_axiClk                                                                      ), //i
    .resetCtrl_axiReset          (resetCtrl_axiReset                                                             )  //i
  );
  Axi4SharedOnChipRam axi_ram (
    .io_axi_arw_valid         (axi_ram_io_axi_arbiter_io_output_arw_valid             ), //i
    .io_axi_arw_ready         (axi_ram_io_axi_arw_ready                               ), //o
    .io_axi_arw_payload_addr  (axi_ram_io_axi_arbiter_io_output_arw_payload_addr[16:0]), //i
    .io_axi_arw_payload_id    (axi_ram_io_axi_arbiter_io_output_arw_payload_id[3:0]   ), //i
    .io_axi_arw_payload_len   (axi_ram_io_axi_arbiter_io_output_arw_payload_len[7:0]  ), //i
    .io_axi_arw_payload_size  (axi_ram_io_axi_arbiter_io_output_arw_payload_size[2:0] ), //i
    .io_axi_arw_payload_burst (axi_ram_io_axi_arbiter_io_output_arw_payload_burst[1:0]), //i
    .io_axi_arw_payload_write (axi_ram_io_axi_arbiter_io_output_arw_payload_write     ), //i
    .io_axi_w_valid           (axi_ram_io_axi_arbiter_io_output_w_valid               ), //i
    .io_axi_w_ready           (axi_ram_io_axi_w_ready                                 ), //o
    .io_axi_w_payload_data    (axi_ram_io_axi_arbiter_io_output_w_payload_data[63:0]  ), //i
    .io_axi_w_payload_strb    (axi_ram_io_axi_arbiter_io_output_w_payload_strb[7:0]   ), //i
    .io_axi_w_payload_last    (axi_ram_io_axi_arbiter_io_output_w_payload_last        ), //i
    .io_axi_b_valid           (axi_ram_io_axi_b_valid                                 ), //o
    .io_axi_b_ready           (axi_ram_io_axi_arbiter_io_output_b_ready               ), //i
    .io_axi_b_payload_id      (axi_ram_io_axi_b_payload_id[3:0]                       ), //o
    .io_axi_b_payload_resp    (axi_ram_io_axi_b_payload_resp[1:0]                     ), //o
    .io_axi_r_valid           (axi_ram_io_axi_r_valid                                 ), //o
    .io_axi_r_ready           (axi_ram_io_axi_arbiter_io_output_r_ready               ), //i
    .io_axi_r_payload_data    (axi_ram_io_axi_r_payload_data[63:0]                    ), //o
    .io_axi_r_payload_id      (axi_ram_io_axi_r_payload_id[3:0]                       ), //o
    .io_axi_r_payload_resp    (axi_ram_io_axi_r_payload_resp[1:0]                     ), //o
    .io_axi_r_payload_last    (axi_ram_io_axi_r_payload_last                          ), //o
    .io_axiClk                (io_axiClk                                              ), //i
    .resetCtrl_axiReset       (resetCtrl_axiReset                                     )  //i
  );
  Axi4SharedOnChipRam_1 axi_bootram (
    .io_axi_arw_valid         (axi_bootram_io_axi_arbiter_io_output_arw_valid             ), //i
    .io_axi_arw_ready         (axi_bootram_io_axi_arw_ready                               ), //o
    .io_axi_arw_payload_addr  (axi_bootram_io_axi_arbiter_io_output_arw_payload_addr[16:0]), //i
    .io_axi_arw_payload_id    (axi_bootram_io_axi_arbiter_io_output_arw_payload_id[3:0]   ), //i
    .io_axi_arw_payload_len   (axi_bootram_io_axi_arbiter_io_output_arw_payload_len[7:0]  ), //i
    .io_axi_arw_payload_size  (axi_bootram_io_axi_arbiter_io_output_arw_payload_size[2:0] ), //i
    .io_axi_arw_payload_burst (axi_bootram_io_axi_arbiter_io_output_arw_payload_burst[1:0]), //i
    .io_axi_arw_payload_write (axi_bootram_io_axi_arbiter_io_output_arw_payload_write     ), //i
    .io_axi_w_valid           (axi_bootram_io_axi_arbiter_io_output_w_valid               ), //i
    .io_axi_w_ready           (axi_bootram_io_axi_w_ready                                 ), //o
    .io_axi_w_payload_data    (axi_bootram_io_axi_arbiter_io_output_w_payload_data[31:0]  ), //i
    .io_axi_w_payload_strb    (axi_bootram_io_axi_arbiter_io_output_w_payload_strb[3:0]   ), //i
    .io_axi_w_payload_last    (axi_bootram_io_axi_arbiter_io_output_w_payload_last        ), //i
    .io_axi_b_valid           (axi_bootram_io_axi_b_valid                                 ), //o
    .io_axi_b_ready           (axi_bootram_io_axi_arbiter_io_output_b_ready               ), //i
    .io_axi_b_payload_id      (axi_bootram_io_axi_b_payload_id[3:0]                       ), //o
    .io_axi_b_payload_resp    (axi_bootram_io_axi_b_payload_resp[1:0]                     ), //o
    .io_axi_r_valid           (axi_bootram_io_axi_r_valid                                 ), //o
    .io_axi_r_ready           (axi_bootram_io_axi_arbiter_io_output_r_ready               ), //i
    .io_axi_r_payload_data    (axi_bootram_io_axi_r_payload_data[31:0]                    ), //o
    .io_axi_r_payload_id      (axi_bootram_io_axi_r_payload_id[3:0]                       ), //o
    .io_axi_r_payload_resp    (axi_bootram_io_axi_r_payload_resp[1:0]                     ), //o
    .io_axi_r_payload_last    (axi_bootram_io_axi_r_payload_last                          ), //o
    .io_axiClk                (io_axiClk                                                  ), //i
    .resetCtrl_axiReset       (resetCtrl_axiReset                                         )  //i
  );
  Axi4SharedToApb3Bridge axi_apbBridge (
    .io_axi_arw_valid         (axi_apbBridge_io_axi_arbiter_io_output_arw_valid             ), //i
    .io_axi_arw_ready         (axi_apbBridge_io_axi_arw_ready                               ), //o
    .io_axi_arw_payload_addr  (axi_apbBridge_io_axi_arbiter_io_output_arw_payload_addr[19:0]), //i
    .io_axi_arw_payload_id    (axi_apbBridge_io_axi_arbiter_io_output_arw_payload_id[3:0]   ), //i
    .io_axi_arw_payload_len   (axi_apbBridge_io_axi_arbiter_io_output_arw_payload_len[7:0]  ), //i
    .io_axi_arw_payload_size  (axi_apbBridge_io_axi_arbiter_io_output_arw_payload_size[2:0] ), //i
    .io_axi_arw_payload_burst (axi_apbBridge_io_axi_arbiter_io_output_arw_payload_burst[1:0]), //i
    .io_axi_arw_payload_write (axi_apbBridge_io_axi_arbiter_io_output_arw_payload_write     ), //i
    .io_axi_w_valid           (axi_apbBridge_io_axi_arbiter_io_output_w_valid               ), //i
    .io_axi_w_ready           (axi_apbBridge_io_axi_w_ready                                 ), //o
    .io_axi_w_payload_data    (axi_apbBridge_io_axi_arbiter_io_output_w_payload_data[31:0]  ), //i
    .io_axi_w_payload_strb    (axi_apbBridge_io_axi_arbiter_io_output_w_payload_strb[3:0]   ), //i
    .io_axi_w_payload_last    (axi_apbBridge_io_axi_arbiter_io_output_w_payload_last        ), //i
    .io_axi_b_valid           (axi_apbBridge_io_axi_b_valid                                 ), //o
    .io_axi_b_ready           (axi_apbBridge_io_axi_arbiter_io_output_b_ready               ), //i
    .io_axi_b_payload_id      (axi_apbBridge_io_axi_b_payload_id[3:0]                       ), //o
    .io_axi_b_payload_resp    (axi_apbBridge_io_axi_b_payload_resp[1:0]                     ), //o
    .io_axi_r_valid           (axi_apbBridge_io_axi_r_valid                                 ), //o
    .io_axi_r_ready           (axi_apbBridge_io_axi_arbiter_io_output_r_ready               ), //i
    .io_axi_r_payload_data    (axi_apbBridge_io_axi_r_payload_data[31:0]                    ), //o
    .io_axi_r_payload_id      (axi_apbBridge_io_axi_r_payload_id[3:0]                       ), //o
    .io_axi_r_payload_resp    (axi_apbBridge_io_axi_r_payload_resp[1:0]                     ), //o
    .io_axi_r_payload_last    (axi_apbBridge_io_axi_r_payload_last                          ), //o
    .io_apb_PADDR             (axi_apbBridge_io_apb_PADDR[19:0]                             ), //o
    .io_apb_PSEL              (axi_apbBridge_io_apb_PSEL                                    ), //o
    .io_apb_PENABLE           (axi_apbBridge_io_apb_PENABLE                                 ), //o
    .io_apb_PREADY            (io_apb_decoder_io_input_PREADY                               ), //i
    .io_apb_PWRITE            (axi_apbBridge_io_apb_PWRITE                                  ), //o
    .io_apb_PWDATA            (axi_apbBridge_io_apb_PWDATA[31:0]                            ), //o
    .io_apb_PRDATA            (io_apb_decoder_io_input_PRDATA[31:0]                         ), //i
    .io_apb_PSLVERROR         (io_apb_decoder_io_input_PSLVERROR                            ), //i
    .io_axiClk                (io_axiClk                                                    ), //i
    .resetCtrl_axiReset       (resetCtrl_axiReset                                           )  //i
  );
  Apb3Uart axi_uartCtrl (
    .io_apb_PADDR     (axi_uartCtrl_io_apb_PADDR[15:0]       ), //i
    .io_apb_PSEL      (apb3Router_1_io_outputs_0_PSEL        ), //i
    .io_apb_PENABLE   (apb3Router_1_io_outputs_0_PENABLE     ), //i
    .io_apb_PREADY    (axi_uartCtrl_io_apb_PREADY            ), //o
    .io_apb_PWRITE    (apb3Router_1_io_outputs_0_PWRITE      ), //i
    .io_apb_PWDATA    (apb3Router_1_io_outputs_0_PWDATA[31:0]), //i
    .io_apb_PRDATA    (axi_uartCtrl_io_apb_PRDATA[31:0]      ), //o
    .io_apb_PSLVERROR (axi_uartCtrl_io_apb_PSLVERROR         ), //o
    .io_uart_txd      (axi_uartCtrl_io_uart_txd              ), //o
    .io_uart_rxd      (io_uart_rxd                           ), //i
    .io_clock         (io_axiClk                             ), //i
    .io_resetn        (axi_uartCtrl_io_resetn                )  //i
  );
  Axi4ReadOnlyDecoder core_cpu_icache_decoder (
    .io_input_ar_valid             (core_cpu_icache_ar_valid                                         ), //i
    .io_input_ar_ready             (core_cpu_icache_decoder_io_input_ar_ready                        ), //o
    .io_input_ar_payload_addr      (core_cpu_icache_ar_payload_addr[63:0]                            ), //i
    .io_input_ar_payload_id        (core_cpu_icache_ar_payload_id[1:0]                               ), //i
    .io_input_ar_payload_len       (core_cpu_icache_ar_payload_len[7:0]                              ), //i
    .io_input_ar_payload_size      (core_cpu_icache_ar_payload_size[2:0]                             ), //i
    .io_input_ar_payload_burst     (core_cpu_icache_ar_payload_burst[1:0]                            ), //i
    .io_input_r_valid              (core_cpu_icache_decoder_io_input_r_valid                         ), //o
    .io_input_r_ready              (core_cpu_icache_r_ready                                          ), //i
    .io_input_r_payload_data       (core_cpu_icache_decoder_io_input_r_payload_data[63:0]            ), //o
    .io_input_r_payload_id         (core_cpu_icache_decoder_io_input_r_payload_id[1:0]               ), //o
    .io_input_r_payload_resp       (core_cpu_icache_decoder_io_input_r_payload_resp[1:0]             ), //o
    .io_input_r_payload_last       (core_cpu_icache_decoder_io_input_r_payload_last                  ), //o
    .io_outputs_0_ar_valid         (core_cpu_icache_decoder_io_outputs_0_ar_valid                    ), //o
    .io_outputs_0_ar_ready         (toplevel_core_cpu_icache_decoder_io_outputs_0_ar_validPipe_fire_1), //i
    .io_outputs_0_ar_payload_addr  (core_cpu_icache_decoder_io_outputs_0_ar_payload_addr[63:0]       ), //o
    .io_outputs_0_ar_payload_id    (core_cpu_icache_decoder_io_outputs_0_ar_payload_id[1:0]          ), //o
    .io_outputs_0_ar_payload_len   (core_cpu_icache_decoder_io_outputs_0_ar_payload_len[7:0]         ), //o
    .io_outputs_0_ar_payload_size  (core_cpu_icache_decoder_io_outputs_0_ar_payload_size[2:0]        ), //o
    .io_outputs_0_ar_payload_burst (core_cpu_icache_decoder_io_outputs_0_ar_payload_burst[1:0]       ), //o
    .io_outputs_0_r_valid          (axi_ram_io_axi_arbiter_io_readInputs_0_r_valid                   ), //i
    .io_outputs_0_r_ready          (core_cpu_icache_decoder_io_outputs_0_r_ready                     ), //o
    .io_outputs_0_r_payload_data   (axi_ram_io_axi_arbiter_io_readInputs_0_r_payload_data[63:0]      ), //i
    .io_outputs_0_r_payload_id     (core_cpu_icache_decoder_io_outputs_0_r_payload_id[1:0]           ), //i
    .io_outputs_0_r_payload_resp   (axi_ram_io_axi_arbiter_io_readInputs_0_r_payload_resp[1:0]       ), //i
    .io_outputs_0_r_payload_last   (axi_ram_io_axi_arbiter_io_readInputs_0_r_payload_last            ), //i
    .io_outputs_1_ar_valid         (core_cpu_icache_decoder_io_outputs_1_ar_valid                    ), //o
    .io_outputs_1_ar_ready         (toplevel_core_cpu_icache_decoder_io_outputs_1_ar_validPipe_fire_1), //i
    .io_outputs_1_ar_payload_addr  (core_cpu_icache_decoder_io_outputs_1_ar_payload_addr[63:0]       ), //o
    .io_outputs_1_ar_payload_id    (core_cpu_icache_decoder_io_outputs_1_ar_payload_id[1:0]          ), //o
    .io_outputs_1_ar_payload_len   (core_cpu_icache_decoder_io_outputs_1_ar_payload_len[7:0]         ), //o
    .io_outputs_1_ar_payload_size  (core_cpu_icache_decoder_io_outputs_1_ar_payload_size[2:0]        ), //o
    .io_outputs_1_ar_payload_burst (core_cpu_icache_decoder_io_outputs_1_ar_payload_burst[1:0]       ), //o
    .io_outputs_1_r_valid          (axi4ReadOnlyArbiter_1_io_inputs_0_r_valid                        ), //i
    .io_outputs_1_r_ready          (core_cpu_icache_decoder_io_outputs_1_r_ready                     ), //o
    .io_outputs_1_r_payload_data   (axi4ReadOnlyArbiter_1_io_inputs_0_r_payload_data[63:0]           ), //i
    .io_outputs_1_r_payload_id     (core_cpu_icache_decoder_io_outputs_1_r_payload_id[1:0]           ), //i
    .io_outputs_1_r_payload_resp   (axi4ReadOnlyArbiter_1_io_inputs_0_r_payload_resp[1:0]            ), //i
    .io_outputs_1_r_payload_last   (axi4ReadOnlyArbiter_1_io_inputs_0_r_payload_last                 ), //i
    .io_axiClk                     (io_axiClk                                                        ), //i
    .resetCtrl_axiReset            (resetCtrl_axiReset                                               )  //i
  );
  Axi4ReadOnlyDecoder core_cpu_dcache_decoder (
    .io_input_ar_valid             (core_cpu_dcache_ar_valid                                         ), //i
    .io_input_ar_ready             (core_cpu_dcache_decoder_io_input_ar_ready                        ), //o
    .io_input_ar_payload_addr      (core_cpu_dcache_ar_payload_addr[63:0]                            ), //i
    .io_input_ar_payload_id        (core_cpu_dcache_ar_payload_id[1:0]                               ), //i
    .io_input_ar_payload_len       (core_cpu_dcache_ar_payload_len[7:0]                              ), //i
    .io_input_ar_payload_size      (core_cpu_dcache_ar_payload_size[2:0]                             ), //i
    .io_input_ar_payload_burst     (core_cpu_dcache_ar_payload_burst[1:0]                            ), //i
    .io_input_r_valid              (core_cpu_dcache_decoder_io_input_r_valid                         ), //o
    .io_input_r_ready              (core_cpu_dcache_r_ready                                          ), //i
    .io_input_r_payload_data       (core_cpu_dcache_decoder_io_input_r_payload_data[63:0]            ), //o
    .io_input_r_payload_id         (core_cpu_dcache_decoder_io_input_r_payload_id[1:0]               ), //o
    .io_input_r_payload_resp       (core_cpu_dcache_decoder_io_input_r_payload_resp[1:0]             ), //o
    .io_input_r_payload_last       (core_cpu_dcache_decoder_io_input_r_payload_last                  ), //o
    .io_outputs_0_ar_valid         (core_cpu_dcache_decoder_io_outputs_0_ar_valid                    ), //o
    .io_outputs_0_ar_ready         (toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_validPipe_fire_1), //i
    .io_outputs_0_ar_payload_addr  (core_cpu_dcache_decoder_io_outputs_0_ar_payload_addr[63:0]       ), //o
    .io_outputs_0_ar_payload_id    (core_cpu_dcache_decoder_io_outputs_0_ar_payload_id[1:0]          ), //o
    .io_outputs_0_ar_payload_len   (core_cpu_dcache_decoder_io_outputs_0_ar_payload_len[7:0]         ), //o
    .io_outputs_0_ar_payload_size  (core_cpu_dcache_decoder_io_outputs_0_ar_payload_size[2:0]        ), //o
    .io_outputs_0_ar_payload_burst (core_cpu_dcache_decoder_io_outputs_0_ar_payload_burst[1:0]       ), //o
    .io_outputs_0_r_valid          (axi_ram_io_axi_arbiter_io_readInputs_1_r_valid                   ), //i
    .io_outputs_0_r_ready          (core_cpu_dcache_decoder_io_outputs_0_r_ready                     ), //o
    .io_outputs_0_r_payload_data   (axi_ram_io_axi_arbiter_io_readInputs_1_r_payload_data[63:0]      ), //i
    .io_outputs_0_r_payload_id     (core_cpu_dcache_decoder_io_outputs_0_r_payload_id[1:0]           ), //i
    .io_outputs_0_r_payload_resp   (axi_ram_io_axi_arbiter_io_readInputs_1_r_payload_resp[1:0]       ), //i
    .io_outputs_0_r_payload_last   (axi_ram_io_axi_arbiter_io_readInputs_1_r_payload_last            ), //i
    .io_outputs_1_ar_valid         (core_cpu_dcache_decoder_io_outputs_1_ar_valid                    ), //o
    .io_outputs_1_ar_ready         (toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_validPipe_fire_1), //i
    .io_outputs_1_ar_payload_addr  (core_cpu_dcache_decoder_io_outputs_1_ar_payload_addr[63:0]       ), //o
    .io_outputs_1_ar_payload_id    (core_cpu_dcache_decoder_io_outputs_1_ar_payload_id[1:0]          ), //o
    .io_outputs_1_ar_payload_len   (core_cpu_dcache_decoder_io_outputs_1_ar_payload_len[7:0]         ), //o
    .io_outputs_1_ar_payload_size  (core_cpu_dcache_decoder_io_outputs_1_ar_payload_size[2:0]        ), //o
    .io_outputs_1_ar_payload_burst (core_cpu_dcache_decoder_io_outputs_1_ar_payload_burst[1:0]       ), //o
    .io_outputs_1_r_valid          (axi4ReadOnlyArbiter_1_io_inputs_1_r_valid                        ), //i
    .io_outputs_1_r_ready          (core_cpu_dcache_decoder_io_outputs_1_r_ready                     ), //o
    .io_outputs_1_r_payload_data   (axi4ReadOnlyArbiter_1_io_inputs_1_r_payload_data[63:0]           ), //i
    .io_outputs_1_r_payload_id     (core_cpu_dcache_decoder_io_outputs_1_r_payload_id[1:0]           ), //i
    .io_outputs_1_r_payload_resp   (axi4ReadOnlyArbiter_1_io_inputs_1_r_payload_resp[1:0]            ), //i
    .io_outputs_1_r_payload_last   (axi4ReadOnlyArbiter_1_io_inputs_1_r_payload_last                 ), //i
    .io_axiClk                     (io_axiClk                                                        ), //i
    .resetCtrl_axiReset            (resetCtrl_axiReset                                               )  //i
  );
  Axi4WriteOnlyDecoder core_cpu_dcache_decoder_1 (
    .io_input_aw_valid             (core_cpu_dcache_aw_valid                                           ), //i
    .io_input_aw_ready             (core_cpu_dcache_decoder_1_io_input_aw_ready                        ), //o
    .io_input_aw_payload_addr      (core_cpu_dcache_aw_payload_addr[63:0]                              ), //i
    .io_input_aw_payload_id        (core_cpu_dcache_aw_payload_id[1:0]                                 ), //i
    .io_input_aw_payload_len       (core_cpu_dcache_aw_payload_len[7:0]                                ), //i
    .io_input_aw_payload_size      (core_cpu_dcache_aw_payload_size[2:0]                               ), //i
    .io_input_aw_payload_burst     (core_cpu_dcache_aw_payload_burst[1:0]                              ), //i
    .io_input_w_valid              (core_cpu_dcache_w_valid                                            ), //i
    .io_input_w_ready              (core_cpu_dcache_decoder_1_io_input_w_ready                         ), //o
    .io_input_w_payload_data       (core_cpu_dcache_w_payload_data[63:0]                               ), //i
    .io_input_w_payload_strb       (core_cpu_dcache_w_payload_strb[7:0]                                ), //i
    .io_input_w_payload_last       (core_cpu_dcache_w_payload_last                                     ), //i
    .io_input_b_valid              (core_cpu_dcache_decoder_1_io_input_b_valid                         ), //o
    .io_input_b_ready              (core_cpu_dcache_b_ready                                            ), //i
    .io_input_b_payload_id         (core_cpu_dcache_decoder_1_io_input_b_payload_id[1:0]               ), //o
    .io_input_b_payload_resp       (core_cpu_dcache_decoder_1_io_input_b_payload_resp[1:0]             ), //o
    .io_outputs_0_aw_valid         (core_cpu_dcache_decoder_1_io_outputs_0_aw_valid                    ), //o
    .io_outputs_0_aw_ready         (toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_validPipe_fire_1), //i
    .io_outputs_0_aw_payload_addr  (core_cpu_dcache_decoder_1_io_outputs_0_aw_payload_addr[63:0]       ), //o
    .io_outputs_0_aw_payload_id    (core_cpu_dcache_decoder_1_io_outputs_0_aw_payload_id[1:0]          ), //o
    .io_outputs_0_aw_payload_len   (core_cpu_dcache_decoder_1_io_outputs_0_aw_payload_len[7:0]         ), //o
    .io_outputs_0_aw_payload_size  (core_cpu_dcache_decoder_1_io_outputs_0_aw_payload_size[2:0]        ), //o
    .io_outputs_0_aw_payload_burst (core_cpu_dcache_decoder_1_io_outputs_0_aw_payload_burst[1:0]       ), //o
    .io_outputs_0_w_valid          (core_cpu_dcache_decoder_1_io_outputs_0_w_valid                     ), //o
    .io_outputs_0_w_ready          (axi_ram_io_axi_arbiter_io_writeInputs_0_w_ready                    ), //i
    .io_outputs_0_w_payload_data   (core_cpu_dcache_decoder_1_io_outputs_0_w_payload_data[63:0]        ), //o
    .io_outputs_0_w_payload_strb   (core_cpu_dcache_decoder_1_io_outputs_0_w_payload_strb[7:0]         ), //o
    .io_outputs_0_w_payload_last   (core_cpu_dcache_decoder_1_io_outputs_0_w_payload_last              ), //o
    .io_outputs_0_b_valid          (axi_ram_io_axi_arbiter_io_writeInputs_0_b_valid                    ), //i
    .io_outputs_0_b_ready          (core_cpu_dcache_decoder_1_io_outputs_0_b_ready                     ), //o
    .io_outputs_0_b_payload_id     (core_cpu_dcache_decoder_1_io_outputs_0_b_payload_id[1:0]           ), //i
    .io_outputs_0_b_payload_resp   (axi_ram_io_axi_arbiter_io_writeInputs_0_b_payload_resp[1:0]        ), //i
    .io_outputs_1_aw_valid         (core_cpu_dcache_decoder_1_io_outputs_1_aw_valid                    ), //o
    .io_outputs_1_aw_ready         (toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_validPipe_fire_1), //i
    .io_outputs_1_aw_payload_addr  (core_cpu_dcache_decoder_1_io_outputs_1_aw_payload_addr[63:0]       ), //o
    .io_outputs_1_aw_payload_id    (core_cpu_dcache_decoder_1_io_outputs_1_aw_payload_id[1:0]          ), //o
    .io_outputs_1_aw_payload_len   (core_cpu_dcache_decoder_1_io_outputs_1_aw_payload_len[7:0]         ), //o
    .io_outputs_1_aw_payload_size  (core_cpu_dcache_decoder_1_io_outputs_1_aw_payload_size[2:0]        ), //o
    .io_outputs_1_aw_payload_burst (core_cpu_dcache_decoder_1_io_outputs_1_aw_payload_burst[1:0]       ), //o
    .io_outputs_1_w_valid          (core_cpu_dcache_decoder_1_io_outputs_1_w_valid                     ), //o
    .io_outputs_1_w_ready          (axi_downsizer_io_input_w_ready                                     ), //i
    .io_outputs_1_w_payload_data   (core_cpu_dcache_decoder_1_io_outputs_1_w_payload_data[63:0]        ), //o
    .io_outputs_1_w_payload_strb   (core_cpu_dcache_decoder_1_io_outputs_1_w_payload_strb[7:0]         ), //o
    .io_outputs_1_w_payload_last   (core_cpu_dcache_decoder_1_io_outputs_1_w_payload_last              ), //o
    .io_outputs_1_b_valid          (axi_downsizer_io_input_b_valid                                     ), //i
    .io_outputs_1_b_ready          (core_cpu_dcache_decoder_1_io_outputs_1_b_ready                     ), //o
    .io_outputs_1_b_payload_id     (core_cpu_dcache_decoder_1_io_outputs_1_b_payload_id[1:0]           ), //i
    .io_outputs_1_b_payload_resp   (axi_downsizer_io_input_b_payload_resp[1:0]                         ), //i
    .io_axiClk                     (io_axiClk                                                          ), //i
    .resetCtrl_axiReset            (resetCtrl_axiReset                                                 )  //i
  );
  Axi4SharedArbiter axi_ram_io_axi_arbiter (
    .io_readInputs_0_ar_valid          (toplevel_core_cpu_icache_decoder_io_outputs_0_ar_validPipe_valid               ), //i
    .io_readInputs_0_ar_ready          (axi_ram_io_axi_arbiter_io_readInputs_0_ar_ready                                ), //o
    .io_readInputs_0_ar_payload_addr   (axi_ram_io_axi_arbiter_io_readInputs_0_ar_payload_addr[16:0]                   ), //i
    .io_readInputs_0_ar_payload_id     (axi_ram_io_axi_arbiter_io_readInputs_0_ar_payload_id[2:0]                      ), //i
    .io_readInputs_0_ar_payload_len    (toplevel_core_cpu_icache_decoder_io_outputs_0_ar_validPipe_payload_len[7:0]    ), //i
    .io_readInputs_0_ar_payload_size   (toplevel_core_cpu_icache_decoder_io_outputs_0_ar_validPipe_payload_size[2:0]   ), //i
    .io_readInputs_0_ar_payload_burst  (toplevel_core_cpu_icache_decoder_io_outputs_0_ar_validPipe_payload_burst[1:0]  ), //i
    .io_readInputs_0_r_valid           (axi_ram_io_axi_arbiter_io_readInputs_0_r_valid                                 ), //o
    .io_readInputs_0_r_ready           (core_cpu_icache_decoder_io_outputs_0_r_ready                                   ), //i
    .io_readInputs_0_r_payload_data    (axi_ram_io_axi_arbiter_io_readInputs_0_r_payload_data[63:0]                    ), //o
    .io_readInputs_0_r_payload_id      (axi_ram_io_axi_arbiter_io_readInputs_0_r_payload_id[2:0]                       ), //o
    .io_readInputs_0_r_payload_resp    (axi_ram_io_axi_arbiter_io_readInputs_0_r_payload_resp[1:0]                     ), //o
    .io_readInputs_0_r_payload_last    (axi_ram_io_axi_arbiter_io_readInputs_0_r_payload_last                          ), //o
    .io_readInputs_1_ar_valid          (toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_validPipe_valid               ), //i
    .io_readInputs_1_ar_ready          (axi_ram_io_axi_arbiter_io_readInputs_1_ar_ready                                ), //o
    .io_readInputs_1_ar_payload_addr   (axi_ram_io_axi_arbiter_io_readInputs_1_ar_payload_addr[16:0]                   ), //i
    .io_readInputs_1_ar_payload_id     (axi_ram_io_axi_arbiter_io_readInputs_1_ar_payload_id[2:0]                      ), //i
    .io_readInputs_1_ar_payload_len    (toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_validPipe_payload_len[7:0]    ), //i
    .io_readInputs_1_ar_payload_size   (toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_validPipe_payload_size[2:0]   ), //i
    .io_readInputs_1_ar_payload_burst  (toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_validPipe_payload_burst[1:0]  ), //i
    .io_readInputs_1_r_valid           (axi_ram_io_axi_arbiter_io_readInputs_1_r_valid                                 ), //o
    .io_readInputs_1_r_ready           (core_cpu_dcache_decoder_io_outputs_0_r_ready                                   ), //i
    .io_readInputs_1_r_payload_data    (axi_ram_io_axi_arbiter_io_readInputs_1_r_payload_data[63:0]                    ), //o
    .io_readInputs_1_r_payload_id      (axi_ram_io_axi_arbiter_io_readInputs_1_r_payload_id[2:0]                       ), //o
    .io_readInputs_1_r_payload_resp    (axi_ram_io_axi_arbiter_io_readInputs_1_r_payload_resp[1:0]                     ), //o
    .io_readInputs_1_r_payload_last    (axi_ram_io_axi_arbiter_io_readInputs_1_r_payload_last                          ), //o
    .io_writeInputs_0_aw_valid         (toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_validPipe_valid             ), //i
    .io_writeInputs_0_aw_ready         (axi_ram_io_axi_arbiter_io_writeInputs_0_aw_ready                               ), //o
    .io_writeInputs_0_aw_payload_addr  (axi_ram_io_axi_arbiter_io_writeInputs_0_aw_payload_addr[16:0]                  ), //i
    .io_writeInputs_0_aw_payload_id    (axi_ram_io_axi_arbiter_io_writeInputs_0_aw_payload_id[3:0]                     ), //i
    .io_writeInputs_0_aw_payload_len   (toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_validPipe_payload_len[7:0]  ), //i
    .io_writeInputs_0_aw_payload_size  (toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_validPipe_payload_size[2:0] ), //i
    .io_writeInputs_0_aw_payload_burst (toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_validPipe_payload_burst[1:0]), //i
    .io_writeInputs_0_w_valid          (core_cpu_dcache_decoder_1_io_outputs_0_w_valid                                 ), //i
    .io_writeInputs_0_w_ready          (axi_ram_io_axi_arbiter_io_writeInputs_0_w_ready                                ), //o
    .io_writeInputs_0_w_payload_data   (core_cpu_dcache_decoder_1_io_outputs_0_w_payload_data[63:0]                    ), //i
    .io_writeInputs_0_w_payload_strb   (core_cpu_dcache_decoder_1_io_outputs_0_w_payload_strb[7:0]                     ), //i
    .io_writeInputs_0_w_payload_last   (core_cpu_dcache_decoder_1_io_outputs_0_w_payload_last                          ), //i
    .io_writeInputs_0_b_valid          (axi_ram_io_axi_arbiter_io_writeInputs_0_b_valid                                ), //o
    .io_writeInputs_0_b_ready          (core_cpu_dcache_decoder_1_io_outputs_0_b_ready                                 ), //i
    .io_writeInputs_0_b_payload_id     (axi_ram_io_axi_arbiter_io_writeInputs_0_b_payload_id[3:0]                      ), //o
    .io_writeInputs_0_b_payload_resp   (axi_ram_io_axi_arbiter_io_writeInputs_0_b_payload_resp[1:0]                    ), //o
    .io_output_arw_valid               (axi_ram_io_axi_arbiter_io_output_arw_valid                                     ), //o
    .io_output_arw_ready               (axi_ram_io_axi_arw_ready                                                       ), //i
    .io_output_arw_payload_addr        (axi_ram_io_axi_arbiter_io_output_arw_payload_addr[16:0]                        ), //o
    .io_output_arw_payload_id          (axi_ram_io_axi_arbiter_io_output_arw_payload_id[3:0]                           ), //o
    .io_output_arw_payload_len         (axi_ram_io_axi_arbiter_io_output_arw_payload_len[7:0]                          ), //o
    .io_output_arw_payload_size        (axi_ram_io_axi_arbiter_io_output_arw_payload_size[2:0]                         ), //o
    .io_output_arw_payload_burst       (axi_ram_io_axi_arbiter_io_output_arw_payload_burst[1:0]                        ), //o
    .io_output_arw_payload_write       (axi_ram_io_axi_arbiter_io_output_arw_payload_write                             ), //o
    .io_output_w_valid                 (axi_ram_io_axi_arbiter_io_output_w_valid                                       ), //o
    .io_output_w_ready                 (axi_ram_io_axi_w_ready                                                         ), //i
    .io_output_w_payload_data          (axi_ram_io_axi_arbiter_io_output_w_payload_data[63:0]                          ), //o
    .io_output_w_payload_strb          (axi_ram_io_axi_arbiter_io_output_w_payload_strb[7:0]                           ), //o
    .io_output_w_payload_last          (axi_ram_io_axi_arbiter_io_output_w_payload_last                                ), //o
    .io_output_b_valid                 (axi_ram_io_axi_b_valid                                                         ), //i
    .io_output_b_ready                 (axi_ram_io_axi_arbiter_io_output_b_ready                                       ), //o
    .io_output_b_payload_id            (axi_ram_io_axi_b_payload_id[3:0]                                               ), //i
    .io_output_b_payload_resp          (axi_ram_io_axi_b_payload_resp[1:0]                                             ), //i
    .io_output_r_valid                 (axi_ram_io_axi_r_valid                                                         ), //i
    .io_output_r_ready                 (axi_ram_io_axi_arbiter_io_output_r_ready                                       ), //o
    .io_output_r_payload_data          (axi_ram_io_axi_r_payload_data[63:0]                                            ), //i
    .io_output_r_payload_id            (axi_ram_io_axi_r_payload_id[3:0]                                               ), //i
    .io_output_r_payload_resp          (axi_ram_io_axi_r_payload_resp[1:0]                                             ), //i
    .io_output_r_payload_last          (axi_ram_io_axi_r_payload_last                                                  ), //i
    .io_axiClk                         (io_axiClk                                                                      ), //i
    .resetCtrl_axiReset                (resetCtrl_axiReset                                                             )  //i
  );
  Axi4ReadOnlyArbiter axi4ReadOnlyArbiter_1 (
    .io_inputs_0_ar_valid          (toplevel_core_cpu_icache_decoder_io_outputs_1_ar_validPipe_valid             ), //i
    .io_inputs_0_ar_ready          (axi4ReadOnlyArbiter_1_io_inputs_0_ar_ready                                   ), //o
    .io_inputs_0_ar_payload_addr   (axi4ReadOnlyArbiter_1_io_inputs_0_ar_payload_addr[31:0]                      ), //i
    .io_inputs_0_ar_payload_id     (axi4ReadOnlyArbiter_1_io_inputs_0_ar_payload_id[2:0]                         ), //i
    .io_inputs_0_ar_payload_region (_zz_io_inputs_0_ar_payload_region[3:0]                                       ), //i
    .io_inputs_0_ar_payload_len    (toplevel_core_cpu_icache_decoder_io_outputs_1_ar_validPipe_payload_len[7:0]  ), //i
    .io_inputs_0_ar_payload_size   (toplevel_core_cpu_icache_decoder_io_outputs_1_ar_validPipe_payload_size[2:0] ), //i
    .io_inputs_0_ar_payload_burst  (toplevel_core_cpu_icache_decoder_io_outputs_1_ar_validPipe_payload_burst[1:0]), //i
    .io_inputs_0_ar_payload_lock   (1'b0                                                                         ), //i
    .io_inputs_0_ar_payload_cache  (4'b0000                                                                      ), //i
    .io_inputs_0_ar_payload_qos    (4'b0000                                                                      ), //i
    .io_inputs_0_ar_payload_prot   (3'b010                                                                       ), //i
    .io_inputs_0_r_valid           (axi4ReadOnlyArbiter_1_io_inputs_0_r_valid                                    ), //o
    .io_inputs_0_r_ready           (core_cpu_icache_decoder_io_outputs_1_r_ready                                 ), //i
    .io_inputs_0_r_payload_data    (axi4ReadOnlyArbiter_1_io_inputs_0_r_payload_data[63:0]                       ), //o
    .io_inputs_0_r_payload_id      (axi4ReadOnlyArbiter_1_io_inputs_0_r_payload_id[2:0]                          ), //o
    .io_inputs_0_r_payload_resp    (axi4ReadOnlyArbiter_1_io_inputs_0_r_payload_resp[1:0]                        ), //o
    .io_inputs_0_r_payload_last    (axi4ReadOnlyArbiter_1_io_inputs_0_r_payload_last                             ), //o
    .io_inputs_1_ar_valid          (toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_validPipe_valid             ), //i
    .io_inputs_1_ar_ready          (axi4ReadOnlyArbiter_1_io_inputs_1_ar_ready                                   ), //o
    .io_inputs_1_ar_payload_addr   (axi4ReadOnlyArbiter_1_io_inputs_1_ar_payload_addr[31:0]                      ), //i
    .io_inputs_1_ar_payload_id     (axi4ReadOnlyArbiter_1_io_inputs_1_ar_payload_id[2:0]                         ), //i
    .io_inputs_1_ar_payload_region (_zz_io_inputs_1_ar_payload_region[3:0]                                       ), //i
    .io_inputs_1_ar_payload_len    (toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_validPipe_payload_len[7:0]  ), //i
    .io_inputs_1_ar_payload_size   (toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_validPipe_payload_size[2:0] ), //i
    .io_inputs_1_ar_payload_burst  (toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_validPipe_payload_burst[1:0]), //i
    .io_inputs_1_ar_payload_lock   (1'b0                                                                         ), //i
    .io_inputs_1_ar_payload_cache  (4'b0000                                                                      ), //i
    .io_inputs_1_ar_payload_qos    (4'b0000                                                                      ), //i
    .io_inputs_1_ar_payload_prot   (3'b010                                                                       ), //i
    .io_inputs_1_r_valid           (axi4ReadOnlyArbiter_1_io_inputs_1_r_valid                                    ), //o
    .io_inputs_1_r_ready           (core_cpu_dcache_decoder_io_outputs_1_r_ready                                 ), //i
    .io_inputs_1_r_payload_data    (axi4ReadOnlyArbiter_1_io_inputs_1_r_payload_data[63:0]                       ), //o
    .io_inputs_1_r_payload_id      (axi4ReadOnlyArbiter_1_io_inputs_1_r_payload_id[2:0]                          ), //o
    .io_inputs_1_r_payload_resp    (axi4ReadOnlyArbiter_1_io_inputs_1_r_payload_resp[1:0]                        ), //o
    .io_inputs_1_r_payload_last    (axi4ReadOnlyArbiter_1_io_inputs_1_r_payload_last                             ), //o
    .io_output_ar_valid            (axi4ReadOnlyArbiter_1_io_output_ar_valid                                     ), //o
    .io_output_ar_ready            (axi_downsizer_io_input_ar_ready                                              ), //i
    .io_output_ar_payload_addr     (axi4ReadOnlyArbiter_1_io_output_ar_payload_addr[31:0]                        ), //o
    .io_output_ar_payload_id       (axi4ReadOnlyArbiter_1_io_output_ar_payload_id[3:0]                           ), //o
    .io_output_ar_payload_region   (axi4ReadOnlyArbiter_1_io_output_ar_payload_region[3:0]                       ), //o
    .io_output_ar_payload_len      (axi4ReadOnlyArbiter_1_io_output_ar_payload_len[7:0]                          ), //o
    .io_output_ar_payload_size     (axi4ReadOnlyArbiter_1_io_output_ar_payload_size[2:0]                         ), //o
    .io_output_ar_payload_burst    (axi4ReadOnlyArbiter_1_io_output_ar_payload_burst[1:0]                        ), //o
    .io_output_ar_payload_lock     (axi4ReadOnlyArbiter_1_io_output_ar_payload_lock                              ), //o
    .io_output_ar_payload_cache    (axi4ReadOnlyArbiter_1_io_output_ar_payload_cache[3:0]                        ), //o
    .io_output_ar_payload_qos      (axi4ReadOnlyArbiter_1_io_output_ar_payload_qos[3:0]                          ), //o
    .io_output_ar_payload_prot     (axi4ReadOnlyArbiter_1_io_output_ar_payload_prot[2:0]                         ), //o
    .io_output_r_valid             (axi_downsizer_io_input_r_valid                                               ), //i
    .io_output_r_ready             (axi4ReadOnlyArbiter_1_io_output_r_ready                                      ), //o
    .io_output_r_payload_data      (axi_downsizer_io_input_r_payload_data[63:0]                                  ), //i
    .io_output_r_payload_id        (axi_downsizer_io_input_r_payload_id[3:0]                                     ), //i
    .io_output_r_payload_resp      (axi_downsizer_io_input_r_payload_resp[1:0]                                   ), //i
    .io_output_r_payload_last      (axi_downsizer_io_input_r_payload_last                                        ), //i
    .io_axiClk                     (io_axiClk                                                                    ), //i
    .resetCtrl_axiReset            (resetCtrl_axiReset                                                           )  //i
  );
  Axi4ReadOnlyDecoder_2 toplevel_axi_downsizer_io_output_readOnly_decoder (
    .io_input_ar_valid              (toplevel_axi_downsizer_io_output_readOnly_ar_valid                                         ), //i
    .io_input_ar_ready              (toplevel_axi_downsizer_io_output_readOnly_decoder_io_input_ar_ready                        ), //o
    .io_input_ar_payload_addr       (toplevel_axi_downsizer_io_output_readOnly_ar_payload_addr[31:0]                            ), //i
    .io_input_ar_payload_id         (toplevel_axi_downsizer_io_output_readOnly_ar_payload_id[3:0]                               ), //i
    .io_input_ar_payload_region     (toplevel_axi_downsizer_io_output_readOnly_ar_payload_region[3:0]                           ), //i
    .io_input_ar_payload_len        (toplevel_axi_downsizer_io_output_readOnly_ar_payload_len[7:0]                              ), //i
    .io_input_ar_payload_size       (toplevel_axi_downsizer_io_output_readOnly_ar_payload_size[2:0]                             ), //i
    .io_input_ar_payload_burst      (toplevel_axi_downsizer_io_output_readOnly_ar_payload_burst[1:0]                            ), //i
    .io_input_ar_payload_lock       (toplevel_axi_downsizer_io_output_readOnly_ar_payload_lock                                  ), //i
    .io_input_ar_payload_cache      (toplevel_axi_downsizer_io_output_readOnly_ar_payload_cache[3:0]                            ), //i
    .io_input_ar_payload_qos        (toplevel_axi_downsizer_io_output_readOnly_ar_payload_qos[3:0]                              ), //i
    .io_input_ar_payload_prot       (toplevel_axi_downsizer_io_output_readOnly_ar_payload_prot[2:0]                             ), //i
    .io_input_r_valid               (toplevel_axi_downsizer_io_output_readOnly_decoder_io_input_r_valid                         ), //o
    .io_input_r_ready               (toplevel_axi_downsizer_io_output_readOnly_r_ready                                          ), //i
    .io_input_r_payload_data        (toplevel_axi_downsizer_io_output_readOnly_decoder_io_input_r_payload_data[31:0]            ), //o
    .io_input_r_payload_id          (toplevel_axi_downsizer_io_output_readOnly_decoder_io_input_r_payload_id[3:0]               ), //o
    .io_input_r_payload_resp        (toplevel_axi_downsizer_io_output_readOnly_decoder_io_input_r_payload_resp[1:0]             ), //o
    .io_input_r_payload_last        (toplevel_axi_downsizer_io_output_readOnly_decoder_io_input_r_payload_last                  ), //o
    .io_outputs_0_ar_valid          (toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_valid                    ), //o
    .io_outputs_0_ar_ready          (toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_fire_1), //i
    .io_outputs_0_ar_payload_addr   (toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_payload_addr[31:0]       ), //o
    .io_outputs_0_ar_payload_id     (toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_payload_id[3:0]          ), //o
    .io_outputs_0_ar_payload_region (toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_payload_region[3:0]      ), //o
    .io_outputs_0_ar_payload_len    (toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_payload_len[7:0]         ), //o
    .io_outputs_0_ar_payload_size   (toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_payload_size[2:0]        ), //o
    .io_outputs_0_ar_payload_burst  (toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_payload_burst[1:0]       ), //o
    .io_outputs_0_ar_payload_lock   (toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_payload_lock             ), //o
    .io_outputs_0_ar_payload_cache  (toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_payload_cache[3:0]       ), //o
    .io_outputs_0_ar_payload_qos    (toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_payload_qos[3:0]         ), //o
    .io_outputs_0_ar_payload_prot   (toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_payload_prot[2:0]        ), //o
    .io_outputs_0_r_valid           (axi_bootram_io_axi_arbiter_io_readInputs_0_r_valid                                         ), //i
    .io_outputs_0_r_ready           (toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_r_ready                     ), //o
    .io_outputs_0_r_payload_data    (axi_bootram_io_axi_arbiter_io_readInputs_0_r_payload_data[31:0]                            ), //i
    .io_outputs_0_r_payload_id      (axi_bootram_io_axi_arbiter_io_readInputs_0_r_payload_id[3:0]                               ), //i
    .io_outputs_0_r_payload_resp    (axi_bootram_io_axi_arbiter_io_readInputs_0_r_payload_resp[1:0]                             ), //i
    .io_outputs_0_r_payload_last    (axi_bootram_io_axi_arbiter_io_readInputs_0_r_payload_last                                  ), //i
    .io_outputs_1_ar_valid          (toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_valid                    ), //o
    .io_outputs_1_ar_ready          (toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_fire_1), //i
    .io_outputs_1_ar_payload_addr   (toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_payload_addr[31:0]       ), //o
    .io_outputs_1_ar_payload_id     (toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_payload_id[3:0]          ), //o
    .io_outputs_1_ar_payload_region (toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_payload_region[3:0]      ), //o
    .io_outputs_1_ar_payload_len    (toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_payload_len[7:0]         ), //o
    .io_outputs_1_ar_payload_size   (toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_payload_size[2:0]        ), //o
    .io_outputs_1_ar_payload_burst  (toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_payload_burst[1:0]       ), //o
    .io_outputs_1_ar_payload_lock   (toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_payload_lock             ), //o
    .io_outputs_1_ar_payload_cache  (toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_payload_cache[3:0]       ), //o
    .io_outputs_1_ar_payload_qos    (toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_payload_qos[3:0]         ), //o
    .io_outputs_1_ar_payload_prot   (toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_payload_prot[2:0]        ), //o
    .io_outputs_1_r_valid           (axi_apbBridge_io_axi_arbiter_io_readInputs_0_r_valid                                       ), //i
    .io_outputs_1_r_ready           (toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_r_ready                     ), //o
    .io_outputs_1_r_payload_data    (axi_apbBridge_io_axi_arbiter_io_readInputs_0_r_payload_data[31:0]                          ), //i
    .io_outputs_1_r_payload_id      (axi_apbBridge_io_axi_arbiter_io_readInputs_0_r_payload_id[3:0]                             ), //i
    .io_outputs_1_r_payload_resp    (axi_apbBridge_io_axi_arbiter_io_readInputs_0_r_payload_resp[1:0]                           ), //i
    .io_outputs_1_r_payload_last    (axi_apbBridge_io_axi_arbiter_io_readInputs_0_r_payload_last                                ), //i
    .io_axiClk                      (io_axiClk                                                                                  ), //i
    .resetCtrl_axiReset             (resetCtrl_axiReset                                                                         )  //i
  );
  Axi4WriteOnlyDecoder_1 toplevel_axi_downsizer_io_output_writeOnly_decoder (
    .io_input_aw_valid              (toplevel_axi_downsizer_io_output_writeOnly_aw_valid                                         ), //i
    .io_input_aw_ready              (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_input_aw_ready                        ), //o
    .io_input_aw_payload_addr       (toplevel_axi_downsizer_io_output_writeOnly_aw_payload_addr[31:0]                            ), //i
    .io_input_aw_payload_id         (toplevel_axi_downsizer_io_output_writeOnly_aw_payload_id[3:0]                               ), //i
    .io_input_aw_payload_region     (toplevel_axi_downsizer_io_output_writeOnly_aw_payload_region[3:0]                           ), //i
    .io_input_aw_payload_len        (toplevel_axi_downsizer_io_output_writeOnly_aw_payload_len[7:0]                              ), //i
    .io_input_aw_payload_size       (toplevel_axi_downsizer_io_output_writeOnly_aw_payload_size[2:0]                             ), //i
    .io_input_aw_payload_burst      (toplevel_axi_downsizer_io_output_writeOnly_aw_payload_burst[1:0]                            ), //i
    .io_input_aw_payload_lock       (toplevel_axi_downsizer_io_output_writeOnly_aw_payload_lock                                  ), //i
    .io_input_aw_payload_cache      (toplevel_axi_downsizer_io_output_writeOnly_aw_payload_cache[3:0]                            ), //i
    .io_input_aw_payload_qos        (toplevel_axi_downsizer_io_output_writeOnly_aw_payload_qos[3:0]                              ), //i
    .io_input_aw_payload_prot       (toplevel_axi_downsizer_io_output_writeOnly_aw_payload_prot[2:0]                             ), //i
    .io_input_w_valid               (toplevel_axi_downsizer_io_output_writeOnly_w_valid                                          ), //i
    .io_input_w_ready               (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_input_w_ready                         ), //o
    .io_input_w_payload_data        (toplevel_axi_downsizer_io_output_writeOnly_w_payload_data[31:0]                             ), //i
    .io_input_w_payload_strb        (toplevel_axi_downsizer_io_output_writeOnly_w_payload_strb[3:0]                              ), //i
    .io_input_w_payload_last        (toplevel_axi_downsizer_io_output_writeOnly_w_payload_last                                   ), //i
    .io_input_b_valid               (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_input_b_valid                         ), //o
    .io_input_b_ready               (toplevel_axi_downsizer_io_output_writeOnly_b_ready                                          ), //i
    .io_input_b_payload_id          (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_input_b_payload_id[3:0]               ), //o
    .io_input_b_payload_resp        (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_input_b_payload_resp[1:0]             ), //o
    .io_outputs_0_aw_valid          (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_valid                    ), //o
    .io_outputs_0_aw_ready          (toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_fire_1), //i
    .io_outputs_0_aw_payload_addr   (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_payload_addr[31:0]       ), //o
    .io_outputs_0_aw_payload_id     (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_payload_id[3:0]          ), //o
    .io_outputs_0_aw_payload_region (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_payload_region[3:0]      ), //o
    .io_outputs_0_aw_payload_len    (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_payload_len[7:0]         ), //o
    .io_outputs_0_aw_payload_size   (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_payload_size[2:0]        ), //o
    .io_outputs_0_aw_payload_burst  (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_payload_burst[1:0]       ), //o
    .io_outputs_0_aw_payload_lock   (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_payload_lock             ), //o
    .io_outputs_0_aw_payload_cache  (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_payload_cache[3:0]       ), //o
    .io_outputs_0_aw_payload_qos    (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_payload_qos[3:0]         ), //o
    .io_outputs_0_aw_payload_prot   (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_payload_prot[2:0]        ), //o
    .io_outputs_0_w_valid           (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_w_valid                     ), //o
    .io_outputs_0_w_ready           (axi_bootram_io_axi_arbiter_io_writeInputs_0_w_ready                                         ), //i
    .io_outputs_0_w_payload_data    (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_w_payload_data[31:0]        ), //o
    .io_outputs_0_w_payload_strb    (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_w_payload_strb[3:0]         ), //o
    .io_outputs_0_w_payload_last    (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_w_payload_last              ), //o
    .io_outputs_0_b_valid           (axi_bootram_io_axi_arbiter_io_writeInputs_0_b_valid                                         ), //i
    .io_outputs_0_b_ready           (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_b_ready                     ), //o
    .io_outputs_0_b_payload_id      (axi_bootram_io_axi_arbiter_io_writeInputs_0_b_payload_id[3:0]                               ), //i
    .io_outputs_0_b_payload_resp    (axi_bootram_io_axi_arbiter_io_writeInputs_0_b_payload_resp[1:0]                             ), //i
    .io_outputs_1_aw_valid          (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_valid                    ), //o
    .io_outputs_1_aw_ready          (toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_fire_1), //i
    .io_outputs_1_aw_payload_addr   (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_payload_addr[31:0]       ), //o
    .io_outputs_1_aw_payload_id     (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_payload_id[3:0]          ), //o
    .io_outputs_1_aw_payload_region (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_payload_region[3:0]      ), //o
    .io_outputs_1_aw_payload_len    (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_payload_len[7:0]         ), //o
    .io_outputs_1_aw_payload_size   (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_payload_size[2:0]        ), //o
    .io_outputs_1_aw_payload_burst  (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_payload_burst[1:0]       ), //o
    .io_outputs_1_aw_payload_lock   (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_payload_lock             ), //o
    .io_outputs_1_aw_payload_cache  (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_payload_cache[3:0]       ), //o
    .io_outputs_1_aw_payload_qos    (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_payload_qos[3:0]         ), //o
    .io_outputs_1_aw_payload_prot   (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_payload_prot[2:0]        ), //o
    .io_outputs_1_w_valid           (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_w_valid                     ), //o
    .io_outputs_1_w_ready           (axi_apbBridge_io_axi_arbiter_io_writeInputs_0_w_ready                                       ), //i
    .io_outputs_1_w_payload_data    (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_w_payload_data[31:0]        ), //o
    .io_outputs_1_w_payload_strb    (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_w_payload_strb[3:0]         ), //o
    .io_outputs_1_w_payload_last    (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_w_payload_last              ), //o
    .io_outputs_1_b_valid           (axi_apbBridge_io_axi_arbiter_io_writeInputs_0_b_valid                                       ), //i
    .io_outputs_1_b_ready           (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_b_ready                     ), //o
    .io_outputs_1_b_payload_id      (axi_apbBridge_io_axi_arbiter_io_writeInputs_0_b_payload_id[3:0]                             ), //i
    .io_outputs_1_b_payload_resp    (axi_apbBridge_io_axi_arbiter_io_writeInputs_0_b_payload_resp[1:0]                           ), //i
    .io_axiClk                      (io_axiClk                                                                                   ), //i
    .resetCtrl_axiReset             (resetCtrl_axiReset                                                                          )  //i
  );
  Axi4SharedArbiter_1 axi_bootram_io_axi_arbiter (
    .io_readInputs_0_ar_valid          (toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_valid              ), //i
    .io_readInputs_0_ar_ready          (axi_bootram_io_axi_arbiter_io_readInputs_0_ar_ready                                                     ), //o
    .io_readInputs_0_ar_payload_addr   (axi_bootram_io_axi_arbiter_io_readInputs_0_ar_payload_addr[16:0]                                        ), //i
    .io_readInputs_0_ar_payload_id     (toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_payload_id[3:0]    ), //i
    .io_readInputs_0_ar_payload_len    (toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_payload_len[7:0]   ), //i
    .io_readInputs_0_ar_payload_size   (toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_payload_size[2:0]  ), //i
    .io_readInputs_0_ar_payload_burst  (toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_payload_burst[1:0] ), //i
    .io_readInputs_0_r_valid           (axi_bootram_io_axi_arbiter_io_readInputs_0_r_valid                                                      ), //o
    .io_readInputs_0_r_ready           (toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_r_ready                                  ), //i
    .io_readInputs_0_r_payload_data    (axi_bootram_io_axi_arbiter_io_readInputs_0_r_payload_data[31:0]                                         ), //o
    .io_readInputs_0_r_payload_id      (axi_bootram_io_axi_arbiter_io_readInputs_0_r_payload_id[3:0]                                            ), //o
    .io_readInputs_0_r_payload_resp    (axi_bootram_io_axi_arbiter_io_readInputs_0_r_payload_resp[1:0]                                          ), //o
    .io_readInputs_0_r_payload_last    (axi_bootram_io_axi_arbiter_io_readInputs_0_r_payload_last                                               ), //o
    .io_writeInputs_0_aw_valid         (toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_valid             ), //i
    .io_writeInputs_0_aw_ready         (axi_bootram_io_axi_arbiter_io_writeInputs_0_aw_ready                                                    ), //o
    .io_writeInputs_0_aw_payload_addr  (axi_bootram_io_axi_arbiter_io_writeInputs_0_aw_payload_addr[16:0]                                       ), //i
    .io_writeInputs_0_aw_payload_id    (toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_id[3:0]   ), //i
    .io_writeInputs_0_aw_payload_len   (toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_len[7:0]  ), //i
    .io_writeInputs_0_aw_payload_size  (toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_size[2:0] ), //i
    .io_writeInputs_0_aw_payload_burst (toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_burst[1:0]), //i
    .io_writeInputs_0_w_valid          (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_w_valid                                 ), //i
    .io_writeInputs_0_w_ready          (axi_bootram_io_axi_arbiter_io_writeInputs_0_w_ready                                                     ), //o
    .io_writeInputs_0_w_payload_data   (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_w_payload_data[31:0]                    ), //i
    .io_writeInputs_0_w_payload_strb   (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_w_payload_strb[3:0]                     ), //i
    .io_writeInputs_0_w_payload_last   (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_w_payload_last                          ), //i
    .io_writeInputs_0_b_valid          (axi_bootram_io_axi_arbiter_io_writeInputs_0_b_valid                                                     ), //o
    .io_writeInputs_0_b_ready          (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_b_ready                                 ), //i
    .io_writeInputs_0_b_payload_id     (axi_bootram_io_axi_arbiter_io_writeInputs_0_b_payload_id[3:0]                                           ), //o
    .io_writeInputs_0_b_payload_resp   (axi_bootram_io_axi_arbiter_io_writeInputs_0_b_payload_resp[1:0]                                         ), //o
    .io_output_arw_valid               (axi_bootram_io_axi_arbiter_io_output_arw_valid                                                          ), //o
    .io_output_arw_ready               (axi_bootram_io_axi_arw_ready                                                                            ), //i
    .io_output_arw_payload_addr        (axi_bootram_io_axi_arbiter_io_output_arw_payload_addr[16:0]                                             ), //o
    .io_output_arw_payload_id          (axi_bootram_io_axi_arbiter_io_output_arw_payload_id[3:0]                                                ), //o
    .io_output_arw_payload_len         (axi_bootram_io_axi_arbiter_io_output_arw_payload_len[7:0]                                               ), //o
    .io_output_arw_payload_size        (axi_bootram_io_axi_arbiter_io_output_arw_payload_size[2:0]                                              ), //o
    .io_output_arw_payload_burst       (axi_bootram_io_axi_arbiter_io_output_arw_payload_burst[1:0]                                             ), //o
    .io_output_arw_payload_write       (axi_bootram_io_axi_arbiter_io_output_arw_payload_write                                                  ), //o
    .io_output_w_valid                 (axi_bootram_io_axi_arbiter_io_output_w_valid                                                            ), //o
    .io_output_w_ready                 (axi_bootram_io_axi_w_ready                                                                              ), //i
    .io_output_w_payload_data          (axi_bootram_io_axi_arbiter_io_output_w_payload_data[31:0]                                               ), //o
    .io_output_w_payload_strb          (axi_bootram_io_axi_arbiter_io_output_w_payload_strb[3:0]                                                ), //o
    .io_output_w_payload_last          (axi_bootram_io_axi_arbiter_io_output_w_payload_last                                                     ), //o
    .io_output_b_valid                 (axi_bootram_io_axi_b_valid                                                                              ), //i
    .io_output_b_ready                 (axi_bootram_io_axi_arbiter_io_output_b_ready                                                            ), //o
    .io_output_b_payload_id            (axi_bootram_io_axi_b_payload_id[3:0]                                                                    ), //i
    .io_output_b_payload_resp          (axi_bootram_io_axi_b_payload_resp[1:0]                                                                  ), //i
    .io_output_r_valid                 (axi_bootram_io_axi_r_valid                                                                              ), //i
    .io_output_r_ready                 (axi_bootram_io_axi_arbiter_io_output_r_ready                                                            ), //o
    .io_output_r_payload_data          (axi_bootram_io_axi_r_payload_data[31:0]                                                                 ), //i
    .io_output_r_payload_id            (axi_bootram_io_axi_r_payload_id[3:0]                                                                    ), //i
    .io_output_r_payload_resp          (axi_bootram_io_axi_r_payload_resp[1:0]                                                                  ), //i
    .io_output_r_payload_last          (axi_bootram_io_axi_r_payload_last                                                                       ), //i
    .io_axiClk                         (io_axiClk                                                                                               ), //i
    .resetCtrl_axiReset                (resetCtrl_axiReset                                                                                      )  //i
  );
  Axi4SharedArbiter_2 axi_apbBridge_io_axi_arbiter (
    .io_readInputs_0_ar_valid          (toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_valid              ), //i
    .io_readInputs_0_ar_ready          (axi_apbBridge_io_axi_arbiter_io_readInputs_0_ar_ready                                                   ), //o
    .io_readInputs_0_ar_payload_addr   (axi_apbBridge_io_axi_arbiter_io_readInputs_0_ar_payload_addr[19:0]                                      ), //i
    .io_readInputs_0_ar_payload_id     (toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_payload_id[3:0]    ), //i
    .io_readInputs_0_ar_payload_len    (toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_payload_len[7:0]   ), //i
    .io_readInputs_0_ar_payload_size   (toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_payload_size[2:0]  ), //i
    .io_readInputs_0_ar_payload_burst  (toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_payload_burst[1:0] ), //i
    .io_readInputs_0_r_valid           (axi_apbBridge_io_axi_arbiter_io_readInputs_0_r_valid                                                    ), //o
    .io_readInputs_0_r_ready           (toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_r_ready                                  ), //i
    .io_readInputs_0_r_payload_data    (axi_apbBridge_io_axi_arbiter_io_readInputs_0_r_payload_data[31:0]                                       ), //o
    .io_readInputs_0_r_payload_id      (axi_apbBridge_io_axi_arbiter_io_readInputs_0_r_payload_id[3:0]                                          ), //o
    .io_readInputs_0_r_payload_resp    (axi_apbBridge_io_axi_arbiter_io_readInputs_0_r_payload_resp[1:0]                                        ), //o
    .io_readInputs_0_r_payload_last    (axi_apbBridge_io_axi_arbiter_io_readInputs_0_r_payload_last                                             ), //o
    .io_writeInputs_0_aw_valid         (toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_valid             ), //i
    .io_writeInputs_0_aw_ready         (axi_apbBridge_io_axi_arbiter_io_writeInputs_0_aw_ready                                                  ), //o
    .io_writeInputs_0_aw_payload_addr  (axi_apbBridge_io_axi_arbiter_io_writeInputs_0_aw_payload_addr[19:0]                                     ), //i
    .io_writeInputs_0_aw_payload_id    (toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_payload_id[3:0]   ), //i
    .io_writeInputs_0_aw_payload_len   (toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_payload_len[7:0]  ), //i
    .io_writeInputs_0_aw_payload_size  (toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_payload_size[2:0] ), //i
    .io_writeInputs_0_aw_payload_burst (toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_payload_burst[1:0]), //i
    .io_writeInputs_0_w_valid          (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_w_valid                                 ), //i
    .io_writeInputs_0_w_ready          (axi_apbBridge_io_axi_arbiter_io_writeInputs_0_w_ready                                                   ), //o
    .io_writeInputs_0_w_payload_data   (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_w_payload_data[31:0]                    ), //i
    .io_writeInputs_0_w_payload_strb   (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_w_payload_strb[3:0]                     ), //i
    .io_writeInputs_0_w_payload_last   (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_w_payload_last                          ), //i
    .io_writeInputs_0_b_valid          (axi_apbBridge_io_axi_arbiter_io_writeInputs_0_b_valid                                                   ), //o
    .io_writeInputs_0_b_ready          (toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_b_ready                                 ), //i
    .io_writeInputs_0_b_payload_id     (axi_apbBridge_io_axi_arbiter_io_writeInputs_0_b_payload_id[3:0]                                         ), //o
    .io_writeInputs_0_b_payload_resp   (axi_apbBridge_io_axi_arbiter_io_writeInputs_0_b_payload_resp[1:0]                                       ), //o
    .io_output_arw_valid               (axi_apbBridge_io_axi_arbiter_io_output_arw_valid                                                        ), //o
    .io_output_arw_ready               (axi_apbBridge_io_axi_arw_ready                                                                          ), //i
    .io_output_arw_payload_addr        (axi_apbBridge_io_axi_arbiter_io_output_arw_payload_addr[19:0]                                           ), //o
    .io_output_arw_payload_id          (axi_apbBridge_io_axi_arbiter_io_output_arw_payload_id[3:0]                                              ), //o
    .io_output_arw_payload_len         (axi_apbBridge_io_axi_arbiter_io_output_arw_payload_len[7:0]                                             ), //o
    .io_output_arw_payload_size        (axi_apbBridge_io_axi_arbiter_io_output_arw_payload_size[2:0]                                            ), //o
    .io_output_arw_payload_burst       (axi_apbBridge_io_axi_arbiter_io_output_arw_payload_burst[1:0]                                           ), //o
    .io_output_arw_payload_write       (axi_apbBridge_io_axi_arbiter_io_output_arw_payload_write                                                ), //o
    .io_output_w_valid                 (axi_apbBridge_io_axi_arbiter_io_output_w_valid                                                          ), //o
    .io_output_w_ready                 (axi_apbBridge_io_axi_w_ready                                                                            ), //i
    .io_output_w_payload_data          (axi_apbBridge_io_axi_arbiter_io_output_w_payload_data[31:0]                                             ), //o
    .io_output_w_payload_strb          (axi_apbBridge_io_axi_arbiter_io_output_w_payload_strb[3:0]                                              ), //o
    .io_output_w_payload_last          (axi_apbBridge_io_axi_arbiter_io_output_w_payload_last                                                   ), //o
    .io_output_b_valid                 (axi_apbBridge_io_axi_b_valid                                                                            ), //i
    .io_output_b_ready                 (axi_apbBridge_io_axi_arbiter_io_output_b_ready                                                          ), //o
    .io_output_b_payload_id            (axi_apbBridge_io_axi_b_payload_id[3:0]                                                                  ), //i
    .io_output_b_payload_resp          (axi_apbBridge_io_axi_b_payload_resp[1:0]                                                                ), //i
    .io_output_r_valid                 (axi_apbBridge_io_axi_r_valid                                                                            ), //i
    .io_output_r_ready                 (axi_apbBridge_io_axi_arbiter_io_output_r_ready                                                          ), //o
    .io_output_r_payload_data          (axi_apbBridge_io_axi_r_payload_data[31:0]                                                               ), //i
    .io_output_r_payload_id            (axi_apbBridge_io_axi_r_payload_id[3:0]                                                                  ), //i
    .io_output_r_payload_resp          (axi_apbBridge_io_axi_r_payload_resp[1:0]                                                                ), //i
    .io_output_r_payload_last          (axi_apbBridge_io_axi_r_payload_last                                                                     ), //i
    .io_axiClk                         (io_axiClk                                                                                               ), //i
    .resetCtrl_axiReset                (resetCtrl_axiReset                                                                                      )  //i
  );
  Apb3Decoder io_apb_decoder (
    .io_input_PADDR      (axi_apbBridge_io_apb_PADDR[19:0]     ), //i
    .io_input_PSEL       (axi_apbBridge_io_apb_PSEL            ), //i
    .io_input_PENABLE    (axi_apbBridge_io_apb_PENABLE         ), //i
    .io_input_PREADY     (io_apb_decoder_io_input_PREADY       ), //o
    .io_input_PWRITE     (axi_apbBridge_io_apb_PWRITE          ), //i
    .io_input_PWDATA     (axi_apbBridge_io_apb_PWDATA[31:0]    ), //i
    .io_input_PRDATA     (io_apb_decoder_io_input_PRDATA[31:0] ), //o
    .io_input_PSLVERROR  (io_apb_decoder_io_input_PSLVERROR    ), //o
    .io_output_PADDR     (io_apb_decoder_io_output_PADDR[19:0] ), //o
    .io_output_PSEL      (io_apb_decoder_io_output_PSEL        ), //o
    .io_output_PENABLE   (io_apb_decoder_io_output_PENABLE     ), //o
    .io_output_PREADY    (apb3Router_1_io_input_PREADY         ), //i
    .io_output_PWRITE    (io_apb_decoder_io_output_PWRITE      ), //o
    .io_output_PWDATA    (io_apb_decoder_io_output_PWDATA[31:0]), //o
    .io_output_PRDATA    (apb3Router_1_io_input_PRDATA[31:0]   ), //i
    .io_output_PSLVERROR (apb3Router_1_io_input_PSLVERROR      )  //i
  );
  Apb3Router apb3Router_1 (
    .io_input_PADDR         (io_apb_decoder_io_output_PADDR[19:0]  ), //i
    .io_input_PSEL          (io_apb_decoder_io_output_PSEL         ), //i
    .io_input_PENABLE       (io_apb_decoder_io_output_PENABLE      ), //i
    .io_input_PREADY        (apb3Router_1_io_input_PREADY          ), //o
    .io_input_PWRITE        (io_apb_decoder_io_output_PWRITE       ), //i
    .io_input_PWDATA        (io_apb_decoder_io_output_PWDATA[31:0] ), //i
    .io_input_PRDATA        (apb3Router_1_io_input_PRDATA[31:0]    ), //o
    .io_input_PSLVERROR     (apb3Router_1_io_input_PSLVERROR       ), //o
    .io_outputs_0_PADDR     (apb3Router_1_io_outputs_0_PADDR[19:0] ), //o
    .io_outputs_0_PSEL      (apb3Router_1_io_outputs_0_PSEL        ), //o
    .io_outputs_0_PENABLE   (apb3Router_1_io_outputs_0_PENABLE     ), //o
    .io_outputs_0_PREADY    (axi_uartCtrl_io_apb_PREADY            ), //i
    .io_outputs_0_PWRITE    (apb3Router_1_io_outputs_0_PWRITE      ), //o
    .io_outputs_0_PWDATA    (apb3Router_1_io_outputs_0_PWDATA[31:0]), //o
    .io_outputs_0_PRDATA    (axi_uartCtrl_io_apb_PRDATA[31:0]      ), //i
    .io_outputs_0_PSLVERROR (axi_uartCtrl_io_apb_PSLVERROR         ), //i
    .io_axiClk              (io_axiClk                             ), //i
    .resetCtrl_axiReset     (resetCtrl_axiReset                    )  //i
  );
  always @(*) begin
    resetCtrl_systemResetUnbuffered = 1'b0;
    if(when_GenDandSocSimple_l89) begin
      resetCtrl_systemResetUnbuffered = 1'b1;
    end
  end

  assign _zz_when_GenDandSocSimple_l89[5 : 0] = 6'h3f;
  assign when_GenDandSocSimple_l89 = (resetCtrl_systemResetCounter != _zz_when_GenDandSocSimple_l89);
  assign bufferCC_1_io_dataIn = (! io_asyncResetn);
  assign when_GenDandSocSimple_l93 = bufferCC_1_io_dataOut;
  assign axi_uartCtrl_io_resetn = (! resetCtrl_axiReset);
  assign axi_downsizer_io_input_aw_payload_addr = toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_validPipe_payload_addr[31:0];
  assign axi_downsizer_io_input_aw_payload_id = {2'd0, toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_validPipe_payload_id};
  assign toplevel_axi_downsizer_io_output_readOnly_ar_valid = axi_downsizer_io_output_ar_valid;
  assign toplevel_axi_downsizer_io_output_readOnly_ar_payload_addr = axi_downsizer_io_output_ar_payload_addr;
  assign toplevel_axi_downsizer_io_output_readOnly_ar_payload_id = axi_downsizer_io_output_ar_payload_id;
  assign toplevel_axi_downsizer_io_output_readOnly_ar_payload_region = axi_downsizer_io_output_ar_payload_region;
  assign toplevel_axi_downsizer_io_output_readOnly_ar_payload_len = axi_downsizer_io_output_ar_payload_len;
  assign toplevel_axi_downsizer_io_output_readOnly_ar_payload_size = axi_downsizer_io_output_ar_payload_size;
  assign toplevel_axi_downsizer_io_output_readOnly_ar_payload_burst = axi_downsizer_io_output_ar_payload_burst;
  assign toplevel_axi_downsizer_io_output_readOnly_ar_payload_lock = axi_downsizer_io_output_ar_payload_lock;
  assign toplevel_axi_downsizer_io_output_readOnly_ar_payload_cache = axi_downsizer_io_output_ar_payload_cache;
  assign toplevel_axi_downsizer_io_output_readOnly_ar_payload_qos = axi_downsizer_io_output_ar_payload_qos;
  assign toplevel_axi_downsizer_io_output_readOnly_ar_payload_prot = axi_downsizer_io_output_ar_payload_prot;
  assign toplevel_axi_downsizer_io_output_readOnly_r_ready = axi_downsizer_io_output_r_ready;
  assign toplevel_axi_downsizer_io_output_writeOnly_aw_valid = axi_downsizer_io_output_aw_valid;
  assign toplevel_axi_downsizer_io_output_writeOnly_aw_payload_addr = axi_downsizer_io_output_aw_payload_addr;
  assign toplevel_axi_downsizer_io_output_writeOnly_aw_payload_id = axi_downsizer_io_output_aw_payload_id;
  assign toplevel_axi_downsizer_io_output_writeOnly_aw_payload_region = axi_downsizer_io_output_aw_payload_region;
  assign toplevel_axi_downsizer_io_output_writeOnly_aw_payload_len = axi_downsizer_io_output_aw_payload_len;
  assign toplevel_axi_downsizer_io_output_writeOnly_aw_payload_size = axi_downsizer_io_output_aw_payload_size;
  assign toplevel_axi_downsizer_io_output_writeOnly_aw_payload_burst = axi_downsizer_io_output_aw_payload_burst;
  assign toplevel_axi_downsizer_io_output_writeOnly_aw_payload_lock = axi_downsizer_io_output_aw_payload_lock;
  assign toplevel_axi_downsizer_io_output_writeOnly_aw_payload_cache = axi_downsizer_io_output_aw_payload_cache;
  assign toplevel_axi_downsizer_io_output_writeOnly_aw_payload_qos = axi_downsizer_io_output_aw_payload_qos;
  assign toplevel_axi_downsizer_io_output_writeOnly_aw_payload_prot = axi_downsizer_io_output_aw_payload_prot;
  assign toplevel_axi_downsizer_io_output_writeOnly_w_valid = axi_downsizer_io_output_w_valid;
  assign toplevel_axi_downsizer_io_output_writeOnly_w_payload_data = axi_downsizer_io_output_w_payload_data;
  assign toplevel_axi_downsizer_io_output_writeOnly_w_payload_strb = axi_downsizer_io_output_w_payload_strb;
  assign toplevel_axi_downsizer_io_output_writeOnly_w_payload_last = axi_downsizer_io_output_w_payload_last;
  assign toplevel_axi_downsizer_io_output_writeOnly_b_ready = axi_downsizer_io_output_b_ready;
  assign toplevel_core_cpu_icache_decoder_io_outputs_0_ar_validPipe_fire = (toplevel_core_cpu_icache_decoder_io_outputs_0_ar_validPipe_valid && toplevel_core_cpu_icache_decoder_io_outputs_0_ar_validPipe_ready);
  assign toplevel_core_cpu_icache_decoder_io_outputs_0_ar_validPipe_fire_1 = (toplevel_core_cpu_icache_decoder_io_outputs_0_ar_validPipe_valid && toplevel_core_cpu_icache_decoder_io_outputs_0_ar_validPipe_ready);
  assign toplevel_core_cpu_icache_decoder_io_outputs_0_ar_validPipe_valid = toplevel_core_cpu_icache_decoder_io_outputs_0_ar_rValid;
  assign toplevel_core_cpu_icache_decoder_io_outputs_0_ar_validPipe_payload_addr = core_cpu_icache_decoder_io_outputs_0_ar_payload_addr;
  assign toplevel_core_cpu_icache_decoder_io_outputs_0_ar_validPipe_payload_id = core_cpu_icache_decoder_io_outputs_0_ar_payload_id;
  assign toplevel_core_cpu_icache_decoder_io_outputs_0_ar_validPipe_payload_len = core_cpu_icache_decoder_io_outputs_0_ar_payload_len;
  assign toplevel_core_cpu_icache_decoder_io_outputs_0_ar_validPipe_payload_size = core_cpu_icache_decoder_io_outputs_0_ar_payload_size;
  assign toplevel_core_cpu_icache_decoder_io_outputs_0_ar_validPipe_payload_burst = core_cpu_icache_decoder_io_outputs_0_ar_payload_burst;
  assign toplevel_core_cpu_icache_decoder_io_outputs_0_ar_validPipe_ready = axi_ram_io_axi_arbiter_io_readInputs_0_ar_ready;
  assign core_cpu_icache_decoder_io_outputs_0_r_payload_id = axi_ram_io_axi_arbiter_io_readInputs_0_r_payload_id[1:0];
  assign toplevel_core_cpu_icache_decoder_io_outputs_1_ar_validPipe_fire = (toplevel_core_cpu_icache_decoder_io_outputs_1_ar_validPipe_valid && toplevel_core_cpu_icache_decoder_io_outputs_1_ar_validPipe_ready);
  assign toplevel_core_cpu_icache_decoder_io_outputs_1_ar_validPipe_fire_1 = (toplevel_core_cpu_icache_decoder_io_outputs_1_ar_validPipe_valid && toplevel_core_cpu_icache_decoder_io_outputs_1_ar_validPipe_ready);
  assign toplevel_core_cpu_icache_decoder_io_outputs_1_ar_validPipe_valid = toplevel_core_cpu_icache_decoder_io_outputs_1_ar_rValid;
  assign toplevel_core_cpu_icache_decoder_io_outputs_1_ar_validPipe_payload_addr = core_cpu_icache_decoder_io_outputs_1_ar_payload_addr;
  assign toplevel_core_cpu_icache_decoder_io_outputs_1_ar_validPipe_payload_id = core_cpu_icache_decoder_io_outputs_1_ar_payload_id;
  assign toplevel_core_cpu_icache_decoder_io_outputs_1_ar_validPipe_payload_len = core_cpu_icache_decoder_io_outputs_1_ar_payload_len;
  assign toplevel_core_cpu_icache_decoder_io_outputs_1_ar_validPipe_payload_size = core_cpu_icache_decoder_io_outputs_1_ar_payload_size;
  assign toplevel_core_cpu_icache_decoder_io_outputs_1_ar_validPipe_payload_burst = core_cpu_icache_decoder_io_outputs_1_ar_payload_burst;
  assign toplevel_core_cpu_icache_decoder_io_outputs_1_ar_validPipe_ready = axi4ReadOnlyArbiter_1_io_inputs_0_ar_ready;
  assign core_cpu_icache_decoder_io_outputs_1_r_payload_id = axi4ReadOnlyArbiter_1_io_inputs_0_r_payload_id[1:0];
  assign toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_validPipe_fire = (toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_validPipe_valid && toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_validPipe_ready);
  assign toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_validPipe_fire_1 = (toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_validPipe_valid && toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_validPipe_ready);
  assign toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_validPipe_valid = toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_rValid;
  assign toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_validPipe_payload_addr = core_cpu_dcache_decoder_io_outputs_0_ar_payload_addr;
  assign toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_validPipe_payload_id = core_cpu_dcache_decoder_io_outputs_0_ar_payload_id;
  assign toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_validPipe_payload_len = core_cpu_dcache_decoder_io_outputs_0_ar_payload_len;
  assign toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_validPipe_payload_size = core_cpu_dcache_decoder_io_outputs_0_ar_payload_size;
  assign toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_validPipe_payload_burst = core_cpu_dcache_decoder_io_outputs_0_ar_payload_burst;
  assign toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_validPipe_ready = axi_ram_io_axi_arbiter_io_readInputs_1_ar_ready;
  assign core_cpu_dcache_decoder_io_outputs_0_r_payload_id = axi_ram_io_axi_arbiter_io_readInputs_1_r_payload_id[1:0];
  assign toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_validPipe_fire = (toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_validPipe_valid && toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_validPipe_ready);
  assign toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_validPipe_fire_1 = (toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_validPipe_valid && toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_validPipe_ready);
  assign toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_validPipe_valid = toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_rValid;
  assign toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_validPipe_payload_addr = core_cpu_dcache_decoder_io_outputs_1_ar_payload_addr;
  assign toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_validPipe_payload_id = core_cpu_dcache_decoder_io_outputs_1_ar_payload_id;
  assign toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_validPipe_payload_len = core_cpu_dcache_decoder_io_outputs_1_ar_payload_len;
  assign toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_validPipe_payload_size = core_cpu_dcache_decoder_io_outputs_1_ar_payload_size;
  assign toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_validPipe_payload_burst = core_cpu_dcache_decoder_io_outputs_1_ar_payload_burst;
  assign toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_validPipe_ready = axi4ReadOnlyArbiter_1_io_inputs_1_ar_ready;
  assign core_cpu_dcache_decoder_io_outputs_1_r_payload_id = axi4ReadOnlyArbiter_1_io_inputs_1_r_payload_id[1:0];
  assign toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_validPipe_fire = (toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_validPipe_valid && toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_validPipe_ready);
  assign toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_validPipe_fire_1 = (toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_validPipe_valid && toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_validPipe_ready);
  assign toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_validPipe_valid = toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_rValid;
  assign toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_validPipe_payload_addr = core_cpu_dcache_decoder_1_io_outputs_0_aw_payload_addr;
  assign toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_validPipe_payload_id = core_cpu_dcache_decoder_1_io_outputs_0_aw_payload_id;
  assign toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_validPipe_payload_len = core_cpu_dcache_decoder_1_io_outputs_0_aw_payload_len;
  assign toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_validPipe_payload_size = core_cpu_dcache_decoder_1_io_outputs_0_aw_payload_size;
  assign toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_validPipe_payload_burst = core_cpu_dcache_decoder_1_io_outputs_0_aw_payload_burst;
  assign toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_validPipe_ready = axi_ram_io_axi_arbiter_io_writeInputs_0_aw_ready;
  assign core_cpu_dcache_decoder_1_io_outputs_0_b_payload_id = axi_ram_io_axi_arbiter_io_writeInputs_0_b_payload_id[1:0];
  assign toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_validPipe_fire = (toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_validPipe_valid && toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_validPipe_ready);
  assign toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_validPipe_fire_1 = (toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_validPipe_valid && toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_validPipe_ready);
  assign toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_validPipe_valid = toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_rValid;
  assign toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_validPipe_payload_addr = core_cpu_dcache_decoder_1_io_outputs_1_aw_payload_addr;
  assign toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_validPipe_payload_id = core_cpu_dcache_decoder_1_io_outputs_1_aw_payload_id;
  assign toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_validPipe_payload_len = core_cpu_dcache_decoder_1_io_outputs_1_aw_payload_len;
  assign toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_validPipe_payload_size = core_cpu_dcache_decoder_1_io_outputs_1_aw_payload_size;
  assign toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_validPipe_payload_burst = core_cpu_dcache_decoder_1_io_outputs_1_aw_payload_burst;
  assign toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_validPipe_ready = axi_downsizer_io_input_aw_ready;
  assign core_cpu_dcache_decoder_1_io_outputs_1_b_payload_id = axi_downsizer_io_input_b_payload_id[1:0];
  assign axi_ram_io_axi_arbiter_io_readInputs_0_ar_payload_addr = toplevel_core_cpu_icache_decoder_io_outputs_0_ar_validPipe_payload_addr[16:0];
  assign axi_ram_io_axi_arbiter_io_readInputs_0_ar_payload_id = {1'd0, toplevel_core_cpu_icache_decoder_io_outputs_0_ar_validPipe_payload_id};
  assign axi_ram_io_axi_arbiter_io_readInputs_1_ar_payload_addr = toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_validPipe_payload_addr[16:0];
  assign axi_ram_io_axi_arbiter_io_readInputs_1_ar_payload_id = {1'd0, toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_validPipe_payload_id};
  assign axi_ram_io_axi_arbiter_io_writeInputs_0_aw_payload_addr = toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_validPipe_payload_addr[16:0];
  assign axi_ram_io_axi_arbiter_io_writeInputs_0_aw_payload_id = {2'd0, toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_validPipe_payload_id};
  assign axi4ReadOnlyArbiter_1_io_inputs_0_ar_payload_addr = toplevel_core_cpu_icache_decoder_io_outputs_1_ar_validPipe_payload_addr[31:0];
  assign axi4ReadOnlyArbiter_1_io_inputs_0_ar_payload_id = {1'd0, toplevel_core_cpu_icache_decoder_io_outputs_1_ar_validPipe_payload_id};
  assign _zz_io_inputs_0_ar_payload_region[3 : 0] = 4'b0000;
  assign axi4ReadOnlyArbiter_1_io_inputs_1_ar_payload_addr = toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_validPipe_payload_addr[31:0];
  assign axi4ReadOnlyArbiter_1_io_inputs_1_ar_payload_id = {1'd0, toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_validPipe_payload_id};
  assign _zz_io_inputs_1_ar_payload_region[3 : 0] = 4'b0000;
  assign _zz_io_input_aw_payload_region[3 : 0] = 4'b0000;
  assign toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_fire = (toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_valid && toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_ready);
  assign toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_fire_1 = (toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_valid && toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_ready);
  assign toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_valid = toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_rValid;
  assign toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_payload_addr = toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_payload_addr;
  assign toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_payload_id = toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_payload_id;
  assign toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_payload_region = toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_payload_region;
  assign toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_payload_len = toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_payload_len;
  assign toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_payload_size = toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_payload_size;
  assign toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_payload_burst = toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_payload_burst;
  assign toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_payload_lock = toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_payload_lock;
  assign toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_payload_cache = toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_payload_cache;
  assign toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_payload_qos = toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_payload_qos;
  assign toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_payload_prot = toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_payload_prot;
  assign toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_ready = axi_bootram_io_axi_arbiter_io_readInputs_0_ar_ready;
  assign toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_fire = (toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_valid && toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_ready);
  assign toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_fire_1 = (toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_valid && toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_ready);
  assign toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_valid = toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_rValid;
  assign toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_payload_addr = toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_payload_addr;
  assign toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_payload_id = toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_payload_id;
  assign toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_payload_region = toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_payload_region;
  assign toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_payload_len = toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_payload_len;
  assign toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_payload_size = toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_payload_size;
  assign toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_payload_burst = toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_payload_burst;
  assign toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_payload_lock = toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_payload_lock;
  assign toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_payload_cache = toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_payload_cache;
  assign toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_payload_qos = toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_payload_qos;
  assign toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_payload_prot = toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_payload_prot;
  assign toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_ready = axi_apbBridge_io_axi_arbiter_io_readInputs_0_ar_ready;
  assign toplevel_axi_downsizer_io_output_readOnly_ar_ready = toplevel_axi_downsizer_io_output_readOnly_decoder_io_input_ar_ready;
  assign toplevel_axi_downsizer_io_output_readOnly_r_valid = toplevel_axi_downsizer_io_output_readOnly_decoder_io_input_r_valid;
  assign toplevel_axi_downsizer_io_output_readOnly_r_payload_data = toplevel_axi_downsizer_io_output_readOnly_decoder_io_input_r_payload_data;
  assign toplevel_axi_downsizer_io_output_readOnly_r_payload_last = toplevel_axi_downsizer_io_output_readOnly_decoder_io_input_r_payload_last;
  assign toplevel_axi_downsizer_io_output_readOnly_r_payload_id = toplevel_axi_downsizer_io_output_readOnly_decoder_io_input_r_payload_id;
  assign toplevel_axi_downsizer_io_output_readOnly_r_payload_resp = toplevel_axi_downsizer_io_output_readOnly_decoder_io_input_r_payload_resp;
  assign toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_fire = (toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_valid && toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_ready);
  assign toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_fire_1 = (toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_valid && toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_ready);
  assign toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_valid = toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_rValid;
  assign toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_addr = toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_payload_addr;
  assign toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_id = toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_payload_id;
  assign toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_region = toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_payload_region;
  assign toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_len = toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_payload_len;
  assign toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_size = toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_payload_size;
  assign toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_burst = toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_payload_burst;
  assign toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_lock = toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_payload_lock;
  assign toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_cache = toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_payload_cache;
  assign toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_qos = toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_payload_qos;
  assign toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_prot = toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_payload_prot;
  assign toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_ready = axi_bootram_io_axi_arbiter_io_writeInputs_0_aw_ready;
  assign toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_fire = (toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_valid && toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_ready);
  assign toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_fire_1 = (toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_valid && toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_ready);
  assign toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_valid = toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_rValid;
  assign toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_payload_addr = toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_payload_addr;
  assign toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_payload_id = toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_payload_id;
  assign toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_payload_region = toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_payload_region;
  assign toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_payload_len = toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_payload_len;
  assign toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_payload_size = toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_payload_size;
  assign toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_payload_burst = toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_payload_burst;
  assign toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_payload_lock = toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_payload_lock;
  assign toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_payload_cache = toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_payload_cache;
  assign toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_payload_qos = toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_payload_qos;
  assign toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_payload_prot = toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_payload_prot;
  assign toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_ready = axi_apbBridge_io_axi_arbiter_io_writeInputs_0_aw_ready;
  assign toplevel_axi_downsizer_io_output_writeOnly_aw_ready = toplevel_axi_downsizer_io_output_writeOnly_decoder_io_input_aw_ready;
  assign toplevel_axi_downsizer_io_output_writeOnly_w_ready = toplevel_axi_downsizer_io_output_writeOnly_decoder_io_input_w_ready;
  assign toplevel_axi_downsizer_io_output_writeOnly_b_valid = toplevel_axi_downsizer_io_output_writeOnly_decoder_io_input_b_valid;
  assign toplevel_axi_downsizer_io_output_writeOnly_b_payload_id = toplevel_axi_downsizer_io_output_writeOnly_decoder_io_input_b_payload_id;
  assign toplevel_axi_downsizer_io_output_writeOnly_b_payload_resp = toplevel_axi_downsizer_io_output_writeOnly_decoder_io_input_b_payload_resp;
  assign axi_bootram_io_axi_arbiter_io_readInputs_0_ar_payload_addr = toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_payload_addr[16:0];
  assign axi_bootram_io_axi_arbiter_io_writeInputs_0_aw_payload_addr = toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_addr[16:0];
  assign axi_apbBridge_io_axi_arbiter_io_readInputs_0_ar_payload_addr = toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_payload_addr[19:0];
  assign axi_apbBridge_io_axi_arbiter_io_writeInputs_0_aw_payload_addr = toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_payload_addr[19:0];
  assign axi_uartCtrl_io_apb_PADDR = apb3Router_1_io_outputs_0_PADDR[15:0];
  assign io_uart_txd = axi_uartCtrl_io_uart_txd;
  always @(posedge io_axiClk or negedge io_asyncResetn) begin
    if(!io_asyncResetn) begin
      resetCtrl_systemResetCounter <= 6'h0;
    end else begin
      if(when_GenDandSocSimple_l89) begin
        resetCtrl_systemResetCounter <= (resetCtrl_systemResetCounter + 6'h01);
      end
      if(when_GenDandSocSimple_l93) begin
        resetCtrl_systemResetCounter <= 6'h0;
      end
    end
  end

  always @(posedge io_axiClk) begin
    resetCtrl_axiReset <= resetCtrl_systemResetUnbuffered;
  end

  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      toplevel_core_cpu_icache_decoder_io_outputs_0_ar_rValid <= 1'b0;
      toplevel_core_cpu_icache_decoder_io_outputs_1_ar_rValid <= 1'b0;
      toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_rValid <= 1'b0;
      toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_rValid <= 1'b0;
      toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_rValid <= 1'b0;
      toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_rValid <= 1'b0;
      toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_rValid <= 1'b0;
      toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_rValid <= 1'b0;
      toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_rValid <= 1'b0;
      toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_rValid <= 1'b0;
    end else begin
      if(core_cpu_icache_decoder_io_outputs_0_ar_valid) begin
        toplevel_core_cpu_icache_decoder_io_outputs_0_ar_rValid <= 1'b1;
      end
      if(toplevel_core_cpu_icache_decoder_io_outputs_0_ar_validPipe_fire) begin
        toplevel_core_cpu_icache_decoder_io_outputs_0_ar_rValid <= 1'b0;
      end
      if(core_cpu_icache_decoder_io_outputs_1_ar_valid) begin
        toplevel_core_cpu_icache_decoder_io_outputs_1_ar_rValid <= 1'b1;
      end
      if(toplevel_core_cpu_icache_decoder_io_outputs_1_ar_validPipe_fire) begin
        toplevel_core_cpu_icache_decoder_io_outputs_1_ar_rValid <= 1'b0;
      end
      if(core_cpu_dcache_decoder_io_outputs_0_ar_valid) begin
        toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_rValid <= 1'b1;
      end
      if(toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_validPipe_fire) begin
        toplevel_core_cpu_dcache_decoder_io_outputs_0_ar_rValid <= 1'b0;
      end
      if(core_cpu_dcache_decoder_io_outputs_1_ar_valid) begin
        toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_rValid <= 1'b1;
      end
      if(toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_validPipe_fire) begin
        toplevel_core_cpu_dcache_decoder_io_outputs_1_ar_rValid <= 1'b0;
      end
      if(core_cpu_dcache_decoder_1_io_outputs_0_aw_valid) begin
        toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_rValid <= 1'b1;
      end
      if(toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_validPipe_fire) begin
        toplevel_core_cpu_dcache_decoder_1_io_outputs_0_aw_rValid <= 1'b0;
      end
      if(core_cpu_dcache_decoder_1_io_outputs_1_aw_valid) begin
        toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_rValid <= 1'b1;
      end
      if(toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_validPipe_fire) begin
        toplevel_core_cpu_dcache_decoder_1_io_outputs_1_aw_rValid <= 1'b0;
      end
      if(toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_valid) begin
        toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_rValid <= 1'b1;
      end
      if(toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_validPipe_fire) begin
        toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_0_ar_rValid <= 1'b0;
      end
      if(toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_valid) begin
        toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_rValid <= 1'b1;
      end
      if(toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_validPipe_fire) begin
        toplevel_toplevel_axi_downsizer_io_output_readOnly_decoder_io_outputs_1_ar_rValid <= 1'b0;
      end
      if(toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_valid) begin
        toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_rValid <= 1'b1;
      end
      if(toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_validPipe_fire) begin
        toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_0_aw_rValid <= 1'b0;
      end
      if(toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_valid) begin
        toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_rValid <= 1'b1;
      end
      if(toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_validPipe_fire) begin
        toplevel_toplevel_axi_downsizer_io_output_writeOnly_decoder_io_outputs_1_aw_rValid <= 1'b0;
      end
    end
  end


endmodule

module Apb3Router (
  input      [19:0]   io_input_PADDR,
  input      [0:0]    io_input_PSEL,
  input               io_input_PENABLE,
  output              io_input_PREADY,
  input               io_input_PWRITE,
  input      [31:0]   io_input_PWDATA,
  output     [31:0]   io_input_PRDATA,
  output              io_input_PSLVERROR,
  output     [19:0]   io_outputs_0_PADDR,
  output     [0:0]    io_outputs_0_PSEL,
  output              io_outputs_0_PENABLE,
  input               io_outputs_0_PREADY,
  output              io_outputs_0_PWRITE,
  output     [31:0]   io_outputs_0_PWDATA,
  input      [31:0]   io_outputs_0_PRDATA,
  input               io_outputs_0_PSLVERROR,
  input               io_axiClk,
  input               resetCtrl_axiReset
);


  assign io_outputs_0_PADDR = io_input_PADDR;
  assign io_outputs_0_PENABLE = io_input_PENABLE;
  assign io_outputs_0_PSEL[0] = io_input_PSEL[0];
  assign io_outputs_0_PWRITE = io_input_PWRITE;
  assign io_outputs_0_PWDATA = io_input_PWDATA;
  assign io_input_PREADY = io_outputs_0_PREADY;
  assign io_input_PRDATA = io_outputs_0_PRDATA;
  assign io_input_PSLVERROR = io_outputs_0_PSLVERROR;

endmodule

module Apb3Decoder (
  input      [19:0]   io_input_PADDR,
  input      [0:0]    io_input_PSEL,
  input               io_input_PENABLE,
  output reg          io_input_PREADY,
  input               io_input_PWRITE,
  input      [31:0]   io_input_PWDATA,
  output     [31:0]   io_input_PRDATA,
  output reg          io_input_PSLVERROR,
  output     [19:0]   io_output_PADDR,
  output     [0:0]    io_output_PSEL,
  output              io_output_PENABLE,
  input               io_output_PREADY,
  output              io_output_PWRITE,
  output     [31:0]   io_output_PWDATA,
  input      [31:0]   io_output_PRDATA,
  input               io_output_PSLVERROR
);

  wire                when_Apb3Decoder_l88;

  assign io_output_PADDR = io_input_PADDR;
  assign io_output_PENABLE = io_input_PENABLE;
  assign io_output_PWRITE = io_input_PWRITE;
  assign io_output_PWDATA = io_input_PWDATA;
  assign io_output_PSEL[0] = (((io_input_PADDR & (~ 20'h00fff)) == 20'h0) && io_input_PSEL[0]);
  always @(*) begin
    io_input_PREADY = io_output_PREADY;
    if(when_Apb3Decoder_l88) begin
      io_input_PREADY = 1'b1;
    end
  end

  assign io_input_PRDATA = io_output_PRDATA;
  always @(*) begin
    io_input_PSLVERROR = io_output_PSLVERROR;
    if(when_Apb3Decoder_l88) begin
      io_input_PSLVERROR = 1'b1;
    end
  end

  assign when_Apb3Decoder_l88 = (io_input_PSEL[0] && (io_output_PSEL == 1'b0));

endmodule

module Axi4SharedArbiter_2 (
  input               io_readInputs_0_ar_valid,
  output              io_readInputs_0_ar_ready,
  input      [19:0]   io_readInputs_0_ar_payload_addr,
  input      [3:0]    io_readInputs_0_ar_payload_id,
  input      [7:0]    io_readInputs_0_ar_payload_len,
  input      [2:0]    io_readInputs_0_ar_payload_size,
  input      [1:0]    io_readInputs_0_ar_payload_burst,
  output              io_readInputs_0_r_valid,
  input               io_readInputs_0_r_ready,
  output     [31:0]   io_readInputs_0_r_payload_data,
  output     [3:0]    io_readInputs_0_r_payload_id,
  output     [1:0]    io_readInputs_0_r_payload_resp,
  output              io_readInputs_0_r_payload_last,
  input               io_writeInputs_0_aw_valid,
  output              io_writeInputs_0_aw_ready,
  input      [19:0]   io_writeInputs_0_aw_payload_addr,
  input      [3:0]    io_writeInputs_0_aw_payload_id,
  input      [7:0]    io_writeInputs_0_aw_payload_len,
  input      [2:0]    io_writeInputs_0_aw_payload_size,
  input      [1:0]    io_writeInputs_0_aw_payload_burst,
  input               io_writeInputs_0_w_valid,
  output              io_writeInputs_0_w_ready,
  input      [31:0]   io_writeInputs_0_w_payload_data,
  input      [3:0]    io_writeInputs_0_w_payload_strb,
  input               io_writeInputs_0_w_payload_last,
  output              io_writeInputs_0_b_valid,
  input               io_writeInputs_0_b_ready,
  output     [3:0]    io_writeInputs_0_b_payload_id,
  output     [1:0]    io_writeInputs_0_b_payload_resp,
  output              io_output_arw_valid,
  input               io_output_arw_ready,
  output     [19:0]   io_output_arw_payload_addr,
  output     [3:0]    io_output_arw_payload_id,
  output     [7:0]    io_output_arw_payload_len,
  output     [2:0]    io_output_arw_payload_size,
  output     [1:0]    io_output_arw_payload_burst,
  output              io_output_arw_payload_write,
  output              io_output_w_valid,
  input               io_output_w_ready,
  output     [31:0]   io_output_w_payload_data,
  output     [3:0]    io_output_w_payload_strb,
  output              io_output_w_payload_last,
  input               io_output_b_valid,
  output              io_output_b_ready,
  input      [3:0]    io_output_b_payload_id,
  input      [1:0]    io_output_b_payload_resp,
  input               io_output_r_valid,
  output              io_output_r_ready,
  input      [31:0]   io_output_r_payload_data,
  input      [3:0]    io_output_r_payload_id,
  input      [1:0]    io_output_r_payload_resp,
  input               io_output_r_payload_last,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  reg                 cmdArbiter_io_output_ready;
  wire                cmdRouteFork_thrown_translated_fifo_io_pop_ready;
  wire                cmdArbiter_io_inputs_0_ready;
  wire                cmdArbiter_io_inputs_1_ready;
  wire                cmdArbiter_io_output_valid;
  wire       [19:0]   cmdArbiter_io_output_payload_addr;
  wire       [3:0]    cmdArbiter_io_output_payload_id;
  wire       [7:0]    cmdArbiter_io_output_payload_len;
  wire       [2:0]    cmdArbiter_io_output_payload_size;
  wire       [1:0]    cmdArbiter_io_output_payload_burst;
  wire                cmdArbiter_io_output_payload_write;
  wire       [0:0]    cmdArbiter_io_chosen;
  wire       [1:0]    cmdArbiter_io_chosenOH;
  wire                cmdRouteFork_thrown_translated_fifo_io_push_ready;
  wire                cmdRouteFork_thrown_translated_fifo_io_pop_valid;
  wire       [2:0]    cmdRouteFork_thrown_translated_fifo_io_occupancy;
  wire                inputsCmd_0_valid;
  wire                inputsCmd_0_ready;
  wire       [19:0]   inputsCmd_0_payload_addr;
  wire       [3:0]    inputsCmd_0_payload_id;
  wire       [7:0]    inputsCmd_0_payload_len;
  wire       [2:0]    inputsCmd_0_payload_size;
  wire       [1:0]    inputsCmd_0_payload_burst;
  wire                inputsCmd_0_payload_write;
  wire                inputsCmd_1_valid;
  wire                inputsCmd_1_ready;
  wire       [19:0]   inputsCmd_1_payload_addr;
  wire       [3:0]    inputsCmd_1_payload_id;
  wire       [7:0]    inputsCmd_1_payload_len;
  wire       [2:0]    inputsCmd_1_payload_size;
  wire       [1:0]    inputsCmd_1_payload_burst;
  wire                inputsCmd_1_payload_write;
  wire                cmdOutputFork_valid;
  wire                cmdOutputFork_ready;
  wire       [19:0]   cmdOutputFork_payload_addr;
  wire       [3:0]    cmdOutputFork_payload_id;
  wire       [7:0]    cmdOutputFork_payload_len;
  wire       [2:0]    cmdOutputFork_payload_size;
  wire       [1:0]    cmdOutputFork_payload_burst;
  wire                cmdOutputFork_payload_write;
  wire                cmdRouteFork_valid;
  reg                 cmdRouteFork_ready;
  wire       [19:0]   cmdRouteFork_payload_addr;
  wire       [3:0]    cmdRouteFork_payload_id;
  wire       [7:0]    cmdRouteFork_payload_len;
  wire       [2:0]    cmdRouteFork_payload_size;
  wire       [1:0]    cmdRouteFork_payload_burst;
  wire                cmdRouteFork_payload_write;
  reg                 axi_apbBridge_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_0;
  reg                 axi_apbBridge_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_1;
  wire                when_Stream_l992;
  wire                when_Stream_l992_1;
  wire                cmdOutputFork_fire;
  wire                cmdRouteFork_fire;
  wire                when_Stream_l438;
  reg                 cmdRouteFork_thrown_valid;
  wire                cmdRouteFork_thrown_ready;
  wire       [19:0]   cmdRouteFork_thrown_payload_addr;
  wire       [3:0]    cmdRouteFork_thrown_payload_id;
  wire       [7:0]    cmdRouteFork_thrown_payload_len;
  wire       [2:0]    cmdRouteFork_thrown_payload_size;
  wire       [1:0]    cmdRouteFork_thrown_payload_burst;
  wire                cmdRouteFork_thrown_payload_write;
  wire                cmdRouteFork_thrown_translated_valid;
  wire                cmdRouteFork_thrown_translated_ready;
  wire                writeLogic_routeDataInput_valid;
  wire                writeLogic_routeDataInput_ready;
  wire       [31:0]   writeLogic_routeDataInput_payload_data;
  wire       [3:0]    writeLogic_routeDataInput_payload_strb;
  wire                writeLogic_routeDataInput_payload_last;
  wire                io_output_w_fire;
  wire                writeLogic_writeRspSels_0;
  wire                readRspSels_0;

  StreamArbiter cmdArbiter (
    .io_inputs_0_valid         (inputsCmd_0_valid                      ), //i
    .io_inputs_0_ready         (cmdArbiter_io_inputs_0_ready           ), //o
    .io_inputs_0_payload_addr  (inputsCmd_0_payload_addr[19:0]         ), //i
    .io_inputs_0_payload_id    (inputsCmd_0_payload_id[3:0]            ), //i
    .io_inputs_0_payload_len   (inputsCmd_0_payload_len[7:0]           ), //i
    .io_inputs_0_payload_size  (inputsCmd_0_payload_size[2:0]          ), //i
    .io_inputs_0_payload_burst (inputsCmd_0_payload_burst[1:0]         ), //i
    .io_inputs_0_payload_write (inputsCmd_0_payload_write              ), //i
    .io_inputs_1_valid         (inputsCmd_1_valid                      ), //i
    .io_inputs_1_ready         (cmdArbiter_io_inputs_1_ready           ), //o
    .io_inputs_1_payload_addr  (inputsCmd_1_payload_addr[19:0]         ), //i
    .io_inputs_1_payload_id    (inputsCmd_1_payload_id[3:0]            ), //i
    .io_inputs_1_payload_len   (inputsCmd_1_payload_len[7:0]           ), //i
    .io_inputs_1_payload_size  (inputsCmd_1_payload_size[2:0]          ), //i
    .io_inputs_1_payload_burst (inputsCmd_1_payload_burst[1:0]         ), //i
    .io_inputs_1_payload_write (inputsCmd_1_payload_write              ), //i
    .io_output_valid           (cmdArbiter_io_output_valid             ), //o
    .io_output_ready           (cmdArbiter_io_output_ready             ), //i
    .io_output_payload_addr    (cmdArbiter_io_output_payload_addr[19:0]), //o
    .io_output_payload_id      (cmdArbiter_io_output_payload_id[3:0]   ), //o
    .io_output_payload_len     (cmdArbiter_io_output_payload_len[7:0]  ), //o
    .io_output_payload_size    (cmdArbiter_io_output_payload_size[2:0] ), //o
    .io_output_payload_burst   (cmdArbiter_io_output_payload_burst[1:0]), //o
    .io_output_payload_write   (cmdArbiter_io_output_payload_write     ), //o
    .io_chosen                 (cmdArbiter_io_chosen                   ), //o
    .io_chosenOH               (cmdArbiter_io_chosenOH[1:0]            ), //o
    .io_axiClk                 (io_axiClk                              ), //i
    .resetCtrl_axiReset        (resetCtrl_axiReset                     )  //i
  );
  StreamFifoLowLatency_2 cmdRouteFork_thrown_translated_fifo (
    .io_push_valid      (cmdRouteFork_thrown_translated_valid                 ), //i
    .io_push_ready      (cmdRouteFork_thrown_translated_fifo_io_push_ready    ), //o
    .io_pop_valid       (cmdRouteFork_thrown_translated_fifo_io_pop_valid     ), //o
    .io_pop_ready       (cmdRouteFork_thrown_translated_fifo_io_pop_ready     ), //i
    .io_flush           (1'b0                                                 ), //i
    .io_occupancy       (cmdRouteFork_thrown_translated_fifo_io_occupancy[2:0]), //o
    .io_axiClk          (io_axiClk                                            ), //i
    .resetCtrl_axiReset (resetCtrl_axiReset                                   )  //i
  );
  assign inputsCmd_0_valid = io_readInputs_0_ar_valid;
  assign io_readInputs_0_ar_ready = inputsCmd_0_ready;
  assign inputsCmd_0_payload_addr = io_readInputs_0_ar_payload_addr;
  assign inputsCmd_0_payload_id = io_readInputs_0_ar_payload_id;
  assign inputsCmd_0_payload_len = io_readInputs_0_ar_payload_len;
  assign inputsCmd_0_payload_size = io_readInputs_0_ar_payload_size;
  assign inputsCmd_0_payload_burst = io_readInputs_0_ar_payload_burst;
  assign inputsCmd_0_payload_write = 1'b0;
  assign inputsCmd_1_valid = io_writeInputs_0_aw_valid;
  assign io_writeInputs_0_aw_ready = inputsCmd_1_ready;
  assign inputsCmd_1_payload_addr = io_writeInputs_0_aw_payload_addr;
  assign inputsCmd_1_payload_id = io_writeInputs_0_aw_payload_id;
  assign inputsCmd_1_payload_len = io_writeInputs_0_aw_payload_len;
  assign inputsCmd_1_payload_size = io_writeInputs_0_aw_payload_size;
  assign inputsCmd_1_payload_burst = io_writeInputs_0_aw_payload_burst;
  assign inputsCmd_1_payload_write = 1'b1;
  assign inputsCmd_0_ready = cmdArbiter_io_inputs_0_ready;
  assign inputsCmd_1_ready = cmdArbiter_io_inputs_1_ready;
  always @(*) begin
    cmdArbiter_io_output_ready = 1'b1;
    if(when_Stream_l992) begin
      cmdArbiter_io_output_ready = 1'b0;
    end
    if(when_Stream_l992_1) begin
      cmdArbiter_io_output_ready = 1'b0;
    end
  end

  assign when_Stream_l992 = ((! cmdOutputFork_ready) && axi_apbBridge_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_0);
  assign when_Stream_l992_1 = ((! cmdRouteFork_ready) && axi_apbBridge_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_1);
  assign cmdOutputFork_valid = (cmdArbiter_io_output_valid && axi_apbBridge_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_0);
  assign cmdOutputFork_payload_addr = cmdArbiter_io_output_payload_addr;
  assign cmdOutputFork_payload_id = cmdArbiter_io_output_payload_id;
  assign cmdOutputFork_payload_len = cmdArbiter_io_output_payload_len;
  assign cmdOutputFork_payload_size = cmdArbiter_io_output_payload_size;
  assign cmdOutputFork_payload_burst = cmdArbiter_io_output_payload_burst;
  assign cmdOutputFork_payload_write = cmdArbiter_io_output_payload_write;
  assign cmdOutputFork_fire = (cmdOutputFork_valid && cmdOutputFork_ready);
  assign cmdRouteFork_valid = (cmdArbiter_io_output_valid && axi_apbBridge_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_1);
  assign cmdRouteFork_payload_addr = cmdArbiter_io_output_payload_addr;
  assign cmdRouteFork_payload_id = cmdArbiter_io_output_payload_id;
  assign cmdRouteFork_payload_len = cmdArbiter_io_output_payload_len;
  assign cmdRouteFork_payload_size = cmdArbiter_io_output_payload_size;
  assign cmdRouteFork_payload_burst = cmdArbiter_io_output_payload_burst;
  assign cmdRouteFork_payload_write = cmdArbiter_io_output_payload_write;
  assign cmdRouteFork_fire = (cmdRouteFork_valid && cmdRouteFork_ready);
  assign io_output_arw_valid = cmdOutputFork_valid;
  assign cmdOutputFork_ready = io_output_arw_ready;
  assign io_output_arw_payload_addr = cmdOutputFork_payload_addr;
  assign io_output_arw_payload_len = cmdOutputFork_payload_len;
  assign io_output_arw_payload_size = cmdOutputFork_payload_size;
  assign io_output_arw_payload_burst = cmdOutputFork_payload_burst;
  assign io_output_arw_payload_write = cmdOutputFork_payload_write;
  assign io_output_arw_payload_id = (cmdOutputFork_payload_write ? cmdOutputFork_payload_id : cmdOutputFork_payload_id);
  assign when_Stream_l438 = (! cmdRouteFork_payload_write);
  always @(*) begin
    cmdRouteFork_thrown_valid = cmdRouteFork_valid;
    if(when_Stream_l438) begin
      cmdRouteFork_thrown_valid = 1'b0;
    end
  end

  always @(*) begin
    cmdRouteFork_ready = cmdRouteFork_thrown_ready;
    if(when_Stream_l438) begin
      cmdRouteFork_ready = 1'b1;
    end
  end

  assign cmdRouteFork_thrown_payload_addr = cmdRouteFork_payload_addr;
  assign cmdRouteFork_thrown_payload_id = cmdRouteFork_payload_id;
  assign cmdRouteFork_thrown_payload_len = cmdRouteFork_payload_len;
  assign cmdRouteFork_thrown_payload_size = cmdRouteFork_payload_size;
  assign cmdRouteFork_thrown_payload_burst = cmdRouteFork_payload_burst;
  assign cmdRouteFork_thrown_payload_write = cmdRouteFork_payload_write;
  assign cmdRouteFork_thrown_translated_valid = cmdRouteFork_thrown_valid;
  assign cmdRouteFork_thrown_ready = cmdRouteFork_thrown_translated_ready;
  assign cmdRouteFork_thrown_translated_ready = cmdRouteFork_thrown_translated_fifo_io_push_ready;
  assign writeLogic_routeDataInput_valid = io_writeInputs_0_w_valid;
  assign writeLogic_routeDataInput_ready = io_writeInputs_0_w_ready;
  assign writeLogic_routeDataInput_payload_data = io_writeInputs_0_w_payload_data;
  assign writeLogic_routeDataInput_payload_strb = io_writeInputs_0_w_payload_strb;
  assign writeLogic_routeDataInput_payload_last = io_writeInputs_0_w_payload_last;
  assign io_output_w_valid = (cmdRouteFork_thrown_translated_fifo_io_pop_valid && writeLogic_routeDataInput_valid);
  assign io_output_w_payload_data = writeLogic_routeDataInput_payload_data;
  assign io_output_w_payload_strb = writeLogic_routeDataInput_payload_strb;
  assign io_output_w_payload_last = writeLogic_routeDataInput_payload_last;
  assign io_writeInputs_0_w_ready = ((cmdRouteFork_thrown_translated_fifo_io_pop_valid && io_output_w_ready) && 1'b1);
  assign io_output_w_fire = (io_output_w_valid && io_output_w_ready);
  assign cmdRouteFork_thrown_translated_fifo_io_pop_ready = (io_output_w_fire && io_output_w_payload_last);
  assign writeLogic_writeRspSels_0 = 1'b1;
  assign io_writeInputs_0_b_valid = (io_output_b_valid && writeLogic_writeRspSels_0);
  assign io_writeInputs_0_b_payload_resp = io_output_b_payload_resp;
  assign io_writeInputs_0_b_payload_id = io_output_b_payload_id;
  assign io_output_b_ready = io_writeInputs_0_b_ready;
  assign readRspSels_0 = 1'b1;
  assign io_readInputs_0_r_valid = (io_output_r_valid && readRspSels_0);
  assign io_readInputs_0_r_payload_data = io_output_r_payload_data;
  assign io_readInputs_0_r_payload_resp = io_output_r_payload_resp;
  assign io_readInputs_0_r_payload_last = io_output_r_payload_last;
  assign io_readInputs_0_r_payload_id = io_output_r_payload_id;
  assign io_output_r_ready = io_readInputs_0_r_ready;
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      axi_apbBridge_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_0 <= 1'b1;
      axi_apbBridge_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_1 <= 1'b1;
    end else begin
      if(cmdOutputFork_fire) begin
        axi_apbBridge_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_0 <= 1'b0;
      end
      if(cmdRouteFork_fire) begin
        axi_apbBridge_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_1 <= 1'b0;
      end
      if(cmdArbiter_io_output_ready) begin
        axi_apbBridge_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_0 <= 1'b1;
        axi_apbBridge_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_1 <= 1'b1;
      end
    end
  end


endmodule

module Axi4SharedArbiter_1 (
  input               io_readInputs_0_ar_valid,
  output              io_readInputs_0_ar_ready,
  input      [16:0]   io_readInputs_0_ar_payload_addr,
  input      [3:0]    io_readInputs_0_ar_payload_id,
  input      [7:0]    io_readInputs_0_ar_payload_len,
  input      [2:0]    io_readInputs_0_ar_payload_size,
  input      [1:0]    io_readInputs_0_ar_payload_burst,
  output              io_readInputs_0_r_valid,
  input               io_readInputs_0_r_ready,
  output     [31:0]   io_readInputs_0_r_payload_data,
  output     [3:0]    io_readInputs_0_r_payload_id,
  output     [1:0]    io_readInputs_0_r_payload_resp,
  output              io_readInputs_0_r_payload_last,
  input               io_writeInputs_0_aw_valid,
  output              io_writeInputs_0_aw_ready,
  input      [16:0]   io_writeInputs_0_aw_payload_addr,
  input      [3:0]    io_writeInputs_0_aw_payload_id,
  input      [7:0]    io_writeInputs_0_aw_payload_len,
  input      [2:0]    io_writeInputs_0_aw_payload_size,
  input      [1:0]    io_writeInputs_0_aw_payload_burst,
  input               io_writeInputs_0_w_valid,
  output              io_writeInputs_0_w_ready,
  input      [31:0]   io_writeInputs_0_w_payload_data,
  input      [3:0]    io_writeInputs_0_w_payload_strb,
  input               io_writeInputs_0_w_payload_last,
  output              io_writeInputs_0_b_valid,
  input               io_writeInputs_0_b_ready,
  output     [3:0]    io_writeInputs_0_b_payload_id,
  output     [1:0]    io_writeInputs_0_b_payload_resp,
  output              io_output_arw_valid,
  input               io_output_arw_ready,
  output     [16:0]   io_output_arw_payload_addr,
  output     [3:0]    io_output_arw_payload_id,
  output     [7:0]    io_output_arw_payload_len,
  output     [2:0]    io_output_arw_payload_size,
  output     [1:0]    io_output_arw_payload_burst,
  output              io_output_arw_payload_write,
  output              io_output_w_valid,
  input               io_output_w_ready,
  output     [31:0]   io_output_w_payload_data,
  output     [3:0]    io_output_w_payload_strb,
  output              io_output_w_payload_last,
  input               io_output_b_valid,
  output              io_output_b_ready,
  input      [3:0]    io_output_b_payload_id,
  input      [1:0]    io_output_b_payload_resp,
  input               io_output_r_valid,
  output              io_output_r_ready,
  input      [31:0]   io_output_r_payload_data,
  input      [3:0]    io_output_r_payload_id,
  input      [1:0]    io_output_r_payload_resp,
  input               io_output_r_payload_last,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  reg                 cmdArbiter_io_output_ready;
  wire                cmdRouteFork_thrown_translated_fifo_io_pop_ready;
  wire                cmdArbiter_io_inputs_0_ready;
  wire                cmdArbiter_io_inputs_1_ready;
  wire                cmdArbiter_io_output_valid;
  wire       [16:0]   cmdArbiter_io_output_payload_addr;
  wire       [3:0]    cmdArbiter_io_output_payload_id;
  wire       [7:0]    cmdArbiter_io_output_payload_len;
  wire       [2:0]    cmdArbiter_io_output_payload_size;
  wire       [1:0]    cmdArbiter_io_output_payload_burst;
  wire                cmdArbiter_io_output_payload_write;
  wire       [0:0]    cmdArbiter_io_chosen;
  wire       [1:0]    cmdArbiter_io_chosenOH;
  wire                cmdRouteFork_thrown_translated_fifo_io_push_ready;
  wire                cmdRouteFork_thrown_translated_fifo_io_pop_valid;
  wire       [2:0]    cmdRouteFork_thrown_translated_fifo_io_occupancy;
  wire                inputsCmd_0_valid;
  wire                inputsCmd_0_ready;
  wire       [16:0]   inputsCmd_0_payload_addr;
  wire       [3:0]    inputsCmd_0_payload_id;
  wire       [7:0]    inputsCmd_0_payload_len;
  wire       [2:0]    inputsCmd_0_payload_size;
  wire       [1:0]    inputsCmd_0_payload_burst;
  wire                inputsCmd_0_payload_write;
  wire                inputsCmd_1_valid;
  wire                inputsCmd_1_ready;
  wire       [16:0]   inputsCmd_1_payload_addr;
  wire       [3:0]    inputsCmd_1_payload_id;
  wire       [7:0]    inputsCmd_1_payload_len;
  wire       [2:0]    inputsCmd_1_payload_size;
  wire       [1:0]    inputsCmd_1_payload_burst;
  wire                inputsCmd_1_payload_write;
  wire                cmdOutputFork_valid;
  wire                cmdOutputFork_ready;
  wire       [16:0]   cmdOutputFork_payload_addr;
  wire       [3:0]    cmdOutputFork_payload_id;
  wire       [7:0]    cmdOutputFork_payload_len;
  wire       [2:0]    cmdOutputFork_payload_size;
  wire       [1:0]    cmdOutputFork_payload_burst;
  wire                cmdOutputFork_payload_write;
  wire                cmdRouteFork_valid;
  reg                 cmdRouteFork_ready;
  wire       [16:0]   cmdRouteFork_payload_addr;
  wire       [3:0]    cmdRouteFork_payload_id;
  wire       [7:0]    cmdRouteFork_payload_len;
  wire       [2:0]    cmdRouteFork_payload_size;
  wire       [1:0]    cmdRouteFork_payload_burst;
  wire                cmdRouteFork_payload_write;
  reg                 axi_bootram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_0;
  reg                 axi_bootram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_1;
  wire                when_Stream_l992;
  wire                when_Stream_l992_1;
  wire                cmdOutputFork_fire;
  wire                cmdRouteFork_fire;
  wire                when_Stream_l438;
  reg                 cmdRouteFork_thrown_valid;
  wire                cmdRouteFork_thrown_ready;
  wire       [16:0]   cmdRouteFork_thrown_payload_addr;
  wire       [3:0]    cmdRouteFork_thrown_payload_id;
  wire       [7:0]    cmdRouteFork_thrown_payload_len;
  wire       [2:0]    cmdRouteFork_thrown_payload_size;
  wire       [1:0]    cmdRouteFork_thrown_payload_burst;
  wire                cmdRouteFork_thrown_payload_write;
  wire                cmdRouteFork_thrown_translated_valid;
  wire                cmdRouteFork_thrown_translated_ready;
  wire                writeLogic_routeDataInput_valid;
  wire                writeLogic_routeDataInput_ready;
  wire       [31:0]   writeLogic_routeDataInput_payload_data;
  wire       [3:0]    writeLogic_routeDataInput_payload_strb;
  wire                writeLogic_routeDataInput_payload_last;
  wire                io_output_w_fire;
  wire                writeLogic_writeRspSels_0;
  wire                readRspSels_0;

  StreamArbiter_1 cmdArbiter (
    .io_inputs_0_valid         (inputsCmd_0_valid                      ), //i
    .io_inputs_0_ready         (cmdArbiter_io_inputs_0_ready           ), //o
    .io_inputs_0_payload_addr  (inputsCmd_0_payload_addr[16:0]         ), //i
    .io_inputs_0_payload_id    (inputsCmd_0_payload_id[3:0]            ), //i
    .io_inputs_0_payload_len   (inputsCmd_0_payload_len[7:0]           ), //i
    .io_inputs_0_payload_size  (inputsCmd_0_payload_size[2:0]          ), //i
    .io_inputs_0_payload_burst (inputsCmd_0_payload_burst[1:0]         ), //i
    .io_inputs_0_payload_write (inputsCmd_0_payload_write              ), //i
    .io_inputs_1_valid         (inputsCmd_1_valid                      ), //i
    .io_inputs_1_ready         (cmdArbiter_io_inputs_1_ready           ), //o
    .io_inputs_1_payload_addr  (inputsCmd_1_payload_addr[16:0]         ), //i
    .io_inputs_1_payload_id    (inputsCmd_1_payload_id[3:0]            ), //i
    .io_inputs_1_payload_len   (inputsCmd_1_payload_len[7:0]           ), //i
    .io_inputs_1_payload_size  (inputsCmd_1_payload_size[2:0]          ), //i
    .io_inputs_1_payload_burst (inputsCmd_1_payload_burst[1:0]         ), //i
    .io_inputs_1_payload_write (inputsCmd_1_payload_write              ), //i
    .io_output_valid           (cmdArbiter_io_output_valid             ), //o
    .io_output_ready           (cmdArbiter_io_output_ready             ), //i
    .io_output_payload_addr    (cmdArbiter_io_output_payload_addr[16:0]), //o
    .io_output_payload_id      (cmdArbiter_io_output_payload_id[3:0]   ), //o
    .io_output_payload_len     (cmdArbiter_io_output_payload_len[7:0]  ), //o
    .io_output_payload_size    (cmdArbiter_io_output_payload_size[2:0] ), //o
    .io_output_payload_burst   (cmdArbiter_io_output_payload_burst[1:0]), //o
    .io_output_payload_write   (cmdArbiter_io_output_payload_write     ), //o
    .io_chosen                 (cmdArbiter_io_chosen                   ), //o
    .io_chosenOH               (cmdArbiter_io_chosenOH[1:0]            ), //o
    .io_axiClk                 (io_axiClk                              ), //i
    .resetCtrl_axiReset        (resetCtrl_axiReset                     )  //i
  );
  StreamFifoLowLatency_2 cmdRouteFork_thrown_translated_fifo (
    .io_push_valid      (cmdRouteFork_thrown_translated_valid                 ), //i
    .io_push_ready      (cmdRouteFork_thrown_translated_fifo_io_push_ready    ), //o
    .io_pop_valid       (cmdRouteFork_thrown_translated_fifo_io_pop_valid     ), //o
    .io_pop_ready       (cmdRouteFork_thrown_translated_fifo_io_pop_ready     ), //i
    .io_flush           (1'b0                                                 ), //i
    .io_occupancy       (cmdRouteFork_thrown_translated_fifo_io_occupancy[2:0]), //o
    .io_axiClk          (io_axiClk                                            ), //i
    .resetCtrl_axiReset (resetCtrl_axiReset                                   )  //i
  );
  assign inputsCmd_0_valid = io_readInputs_0_ar_valid;
  assign io_readInputs_0_ar_ready = inputsCmd_0_ready;
  assign inputsCmd_0_payload_addr = io_readInputs_0_ar_payload_addr;
  assign inputsCmd_0_payload_id = io_readInputs_0_ar_payload_id;
  assign inputsCmd_0_payload_len = io_readInputs_0_ar_payload_len;
  assign inputsCmd_0_payload_size = io_readInputs_0_ar_payload_size;
  assign inputsCmd_0_payload_burst = io_readInputs_0_ar_payload_burst;
  assign inputsCmd_0_payload_write = 1'b0;
  assign inputsCmd_1_valid = io_writeInputs_0_aw_valid;
  assign io_writeInputs_0_aw_ready = inputsCmd_1_ready;
  assign inputsCmd_1_payload_addr = io_writeInputs_0_aw_payload_addr;
  assign inputsCmd_1_payload_id = io_writeInputs_0_aw_payload_id;
  assign inputsCmd_1_payload_len = io_writeInputs_0_aw_payload_len;
  assign inputsCmd_1_payload_size = io_writeInputs_0_aw_payload_size;
  assign inputsCmd_1_payload_burst = io_writeInputs_0_aw_payload_burst;
  assign inputsCmd_1_payload_write = 1'b1;
  assign inputsCmd_0_ready = cmdArbiter_io_inputs_0_ready;
  assign inputsCmd_1_ready = cmdArbiter_io_inputs_1_ready;
  always @(*) begin
    cmdArbiter_io_output_ready = 1'b1;
    if(when_Stream_l992) begin
      cmdArbiter_io_output_ready = 1'b0;
    end
    if(when_Stream_l992_1) begin
      cmdArbiter_io_output_ready = 1'b0;
    end
  end

  assign when_Stream_l992 = ((! cmdOutputFork_ready) && axi_bootram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_0);
  assign when_Stream_l992_1 = ((! cmdRouteFork_ready) && axi_bootram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_1);
  assign cmdOutputFork_valid = (cmdArbiter_io_output_valid && axi_bootram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_0);
  assign cmdOutputFork_payload_addr = cmdArbiter_io_output_payload_addr;
  assign cmdOutputFork_payload_id = cmdArbiter_io_output_payload_id;
  assign cmdOutputFork_payload_len = cmdArbiter_io_output_payload_len;
  assign cmdOutputFork_payload_size = cmdArbiter_io_output_payload_size;
  assign cmdOutputFork_payload_burst = cmdArbiter_io_output_payload_burst;
  assign cmdOutputFork_payload_write = cmdArbiter_io_output_payload_write;
  assign cmdOutputFork_fire = (cmdOutputFork_valid && cmdOutputFork_ready);
  assign cmdRouteFork_valid = (cmdArbiter_io_output_valid && axi_bootram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_1);
  assign cmdRouteFork_payload_addr = cmdArbiter_io_output_payload_addr;
  assign cmdRouteFork_payload_id = cmdArbiter_io_output_payload_id;
  assign cmdRouteFork_payload_len = cmdArbiter_io_output_payload_len;
  assign cmdRouteFork_payload_size = cmdArbiter_io_output_payload_size;
  assign cmdRouteFork_payload_burst = cmdArbiter_io_output_payload_burst;
  assign cmdRouteFork_payload_write = cmdArbiter_io_output_payload_write;
  assign cmdRouteFork_fire = (cmdRouteFork_valid && cmdRouteFork_ready);
  assign io_output_arw_valid = cmdOutputFork_valid;
  assign cmdOutputFork_ready = io_output_arw_ready;
  assign io_output_arw_payload_addr = cmdOutputFork_payload_addr;
  assign io_output_arw_payload_len = cmdOutputFork_payload_len;
  assign io_output_arw_payload_size = cmdOutputFork_payload_size;
  assign io_output_arw_payload_burst = cmdOutputFork_payload_burst;
  assign io_output_arw_payload_write = cmdOutputFork_payload_write;
  assign io_output_arw_payload_id = (cmdOutputFork_payload_write ? cmdOutputFork_payload_id : cmdOutputFork_payload_id);
  assign when_Stream_l438 = (! cmdRouteFork_payload_write);
  always @(*) begin
    cmdRouteFork_thrown_valid = cmdRouteFork_valid;
    if(when_Stream_l438) begin
      cmdRouteFork_thrown_valid = 1'b0;
    end
  end

  always @(*) begin
    cmdRouteFork_ready = cmdRouteFork_thrown_ready;
    if(when_Stream_l438) begin
      cmdRouteFork_ready = 1'b1;
    end
  end

  assign cmdRouteFork_thrown_payload_addr = cmdRouteFork_payload_addr;
  assign cmdRouteFork_thrown_payload_id = cmdRouteFork_payload_id;
  assign cmdRouteFork_thrown_payload_len = cmdRouteFork_payload_len;
  assign cmdRouteFork_thrown_payload_size = cmdRouteFork_payload_size;
  assign cmdRouteFork_thrown_payload_burst = cmdRouteFork_payload_burst;
  assign cmdRouteFork_thrown_payload_write = cmdRouteFork_payload_write;
  assign cmdRouteFork_thrown_translated_valid = cmdRouteFork_thrown_valid;
  assign cmdRouteFork_thrown_ready = cmdRouteFork_thrown_translated_ready;
  assign cmdRouteFork_thrown_translated_ready = cmdRouteFork_thrown_translated_fifo_io_push_ready;
  assign writeLogic_routeDataInput_valid = io_writeInputs_0_w_valid;
  assign writeLogic_routeDataInput_ready = io_writeInputs_0_w_ready;
  assign writeLogic_routeDataInput_payload_data = io_writeInputs_0_w_payload_data;
  assign writeLogic_routeDataInput_payload_strb = io_writeInputs_0_w_payload_strb;
  assign writeLogic_routeDataInput_payload_last = io_writeInputs_0_w_payload_last;
  assign io_output_w_valid = (cmdRouteFork_thrown_translated_fifo_io_pop_valid && writeLogic_routeDataInput_valid);
  assign io_output_w_payload_data = writeLogic_routeDataInput_payload_data;
  assign io_output_w_payload_strb = writeLogic_routeDataInput_payload_strb;
  assign io_output_w_payload_last = writeLogic_routeDataInput_payload_last;
  assign io_writeInputs_0_w_ready = ((cmdRouteFork_thrown_translated_fifo_io_pop_valid && io_output_w_ready) && 1'b1);
  assign io_output_w_fire = (io_output_w_valid && io_output_w_ready);
  assign cmdRouteFork_thrown_translated_fifo_io_pop_ready = (io_output_w_fire && io_output_w_payload_last);
  assign writeLogic_writeRspSels_0 = 1'b1;
  assign io_writeInputs_0_b_valid = (io_output_b_valid && writeLogic_writeRspSels_0);
  assign io_writeInputs_0_b_payload_resp = io_output_b_payload_resp;
  assign io_writeInputs_0_b_payload_id = io_output_b_payload_id;
  assign io_output_b_ready = io_writeInputs_0_b_ready;
  assign readRspSels_0 = 1'b1;
  assign io_readInputs_0_r_valid = (io_output_r_valid && readRspSels_0);
  assign io_readInputs_0_r_payload_data = io_output_r_payload_data;
  assign io_readInputs_0_r_payload_resp = io_output_r_payload_resp;
  assign io_readInputs_0_r_payload_last = io_output_r_payload_last;
  assign io_readInputs_0_r_payload_id = io_output_r_payload_id;
  assign io_output_r_ready = io_readInputs_0_r_ready;
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      axi_bootram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_0 <= 1'b1;
      axi_bootram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_1 <= 1'b1;
    end else begin
      if(cmdOutputFork_fire) begin
        axi_bootram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_0 <= 1'b0;
      end
      if(cmdRouteFork_fire) begin
        axi_bootram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_1 <= 1'b0;
      end
      if(cmdArbiter_io_output_ready) begin
        axi_bootram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_0 <= 1'b1;
        axi_bootram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_1 <= 1'b1;
      end
    end
  end


endmodule

module Axi4WriteOnlyDecoder_1 (
  input               io_input_aw_valid,
  output              io_input_aw_ready,
  input      [31:0]   io_input_aw_payload_addr,
  input      [3:0]    io_input_aw_payload_id,
  input      [3:0]    io_input_aw_payload_region,
  input      [7:0]    io_input_aw_payload_len,
  input      [2:0]    io_input_aw_payload_size,
  input      [1:0]    io_input_aw_payload_burst,
  input      [0:0]    io_input_aw_payload_lock,
  input      [3:0]    io_input_aw_payload_cache,
  input      [3:0]    io_input_aw_payload_qos,
  input      [2:0]    io_input_aw_payload_prot,
  input               io_input_w_valid,
  output              io_input_w_ready,
  input      [31:0]   io_input_w_payload_data,
  input      [3:0]    io_input_w_payload_strb,
  input               io_input_w_payload_last,
  output              io_input_b_valid,
  input               io_input_b_ready,
  output reg [3:0]    io_input_b_payload_id,
  output reg [1:0]    io_input_b_payload_resp,
  output              io_outputs_0_aw_valid,
  input               io_outputs_0_aw_ready,
  output     [31:0]   io_outputs_0_aw_payload_addr,
  output     [3:0]    io_outputs_0_aw_payload_id,
  output     [3:0]    io_outputs_0_aw_payload_region,
  output     [7:0]    io_outputs_0_aw_payload_len,
  output     [2:0]    io_outputs_0_aw_payload_size,
  output     [1:0]    io_outputs_0_aw_payload_burst,
  output     [0:0]    io_outputs_0_aw_payload_lock,
  output     [3:0]    io_outputs_0_aw_payload_cache,
  output     [3:0]    io_outputs_0_aw_payload_qos,
  output     [2:0]    io_outputs_0_aw_payload_prot,
  output              io_outputs_0_w_valid,
  input               io_outputs_0_w_ready,
  output     [31:0]   io_outputs_0_w_payload_data,
  output     [3:0]    io_outputs_0_w_payload_strb,
  output              io_outputs_0_w_payload_last,
  input               io_outputs_0_b_valid,
  output              io_outputs_0_b_ready,
  input      [3:0]    io_outputs_0_b_payload_id,
  input      [1:0]    io_outputs_0_b_payload_resp,
  output              io_outputs_1_aw_valid,
  input               io_outputs_1_aw_ready,
  output     [31:0]   io_outputs_1_aw_payload_addr,
  output     [3:0]    io_outputs_1_aw_payload_id,
  output     [3:0]    io_outputs_1_aw_payload_region,
  output     [7:0]    io_outputs_1_aw_payload_len,
  output     [2:0]    io_outputs_1_aw_payload_size,
  output     [1:0]    io_outputs_1_aw_payload_burst,
  output     [0:0]    io_outputs_1_aw_payload_lock,
  output     [3:0]    io_outputs_1_aw_payload_cache,
  output     [3:0]    io_outputs_1_aw_payload_qos,
  output     [2:0]    io_outputs_1_aw_payload_prot,
  output              io_outputs_1_w_valid,
  input               io_outputs_1_w_ready,
  output     [31:0]   io_outputs_1_w_payload_data,
  output     [3:0]    io_outputs_1_w_payload_strb,
  output              io_outputs_1_w_payload_last,
  input               io_outputs_1_b_valid,
  output              io_outputs_1_b_ready,
  input      [3:0]    io_outputs_1_b_payload_id,
  input      [1:0]    io_outputs_1_b_payload_resp,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  wire                errorSlave_io_axi_aw_valid;
  wire                errorSlave_io_axi_w_valid;
  wire                errorSlave_io_axi_aw_ready;
  wire                errorSlave_io_axi_w_ready;
  wire                errorSlave_io_axi_b_valid;
  wire       [3:0]    errorSlave_io_axi_b_payload_id;
  wire       [1:0]    errorSlave_io_axi_b_payload_resp;
  wire                cmdAllowedStart;
  wire                io_input_aw_fire;
  wire                io_input_b_fire;
  reg                 pendingCmdCounter_incrementIt;
  reg                 pendingCmdCounter_decrementIt;
  wire       [2:0]    pendingCmdCounter_valueNext;
  reg        [2:0]    pendingCmdCounter_value;
  wire                pendingCmdCounter_willOverflowIfInc;
  wire                pendingCmdCounter_willOverflow;
  reg        [2:0]    pendingCmdCounter_finalIncrement;
  wire                when_Utils_l669;
  wire                when_Utils_l671;
  wire                io_input_w_fire;
  wire                when_Utils_l644;
  reg                 pendingDataCounter_incrementIt;
  reg                 pendingDataCounter_decrementIt;
  wire       [2:0]    pendingDataCounter_valueNext;
  reg        [2:0]    pendingDataCounter_value;
  wire                pendingDataCounter_willOverflowIfInc;
  wire                pendingDataCounter_willOverflow;
  reg        [2:0]    pendingDataCounter_finalIncrement;
  wire                when_Utils_l669_1;
  wire                when_Utils_l671_1;
  wire       [1:0]    decodedCmdSels;
  wire                decodedCmdError;
  reg        [1:0]    pendingSels;
  reg                 pendingError;
  wire                allowCmd;
  wire                allowData;
  reg                 _zz_cmdAllowedStart;
  wire                _zz_io_input_b_payload_id;
  wire                _zz_io_outputs_1_w_valid;
  wire       [0:0]    writeRspIndex;

  Axi4WriteOnlyErrorSlave errorSlave (
    .io_axi_aw_valid          (errorSlave_io_axi_aw_valid           ), //i
    .io_axi_aw_ready          (errorSlave_io_axi_aw_ready           ), //o
    .io_axi_aw_payload_addr   (io_input_aw_payload_addr[31:0]       ), //i
    .io_axi_aw_payload_id     (io_input_aw_payload_id[3:0]          ), //i
    .io_axi_aw_payload_region (io_input_aw_payload_region[3:0]      ), //i
    .io_axi_aw_payload_len    (io_input_aw_payload_len[7:0]         ), //i
    .io_axi_aw_payload_size   (io_input_aw_payload_size[2:0]        ), //i
    .io_axi_aw_payload_burst  (io_input_aw_payload_burst[1:0]       ), //i
    .io_axi_aw_payload_lock   (io_input_aw_payload_lock             ), //i
    .io_axi_aw_payload_cache  (io_input_aw_payload_cache[3:0]       ), //i
    .io_axi_aw_payload_qos    (io_input_aw_payload_qos[3:0]         ), //i
    .io_axi_aw_payload_prot   (io_input_aw_payload_prot[2:0]        ), //i
    .io_axi_w_valid           (errorSlave_io_axi_w_valid            ), //i
    .io_axi_w_ready           (errorSlave_io_axi_w_ready            ), //o
    .io_axi_w_payload_data    (io_input_w_payload_data[31:0]        ), //i
    .io_axi_w_payload_strb    (io_input_w_payload_strb[3:0]         ), //i
    .io_axi_w_payload_last    (io_input_w_payload_last              ), //i
    .io_axi_b_valid           (errorSlave_io_axi_b_valid            ), //o
    .io_axi_b_ready           (io_input_b_ready                     ), //i
    .io_axi_b_payload_id      (errorSlave_io_axi_b_payload_id[3:0]  ), //o
    .io_axi_b_payload_resp    (errorSlave_io_axi_b_payload_resp[1:0]), //o
    .io_axiClk                (io_axiClk                            ), //i
    .resetCtrl_axiReset       (resetCtrl_axiReset                   )  //i
  );
  assign io_input_aw_fire = (io_input_aw_valid && io_input_aw_ready);
  assign io_input_b_fire = (io_input_b_valid && io_input_b_ready);
  always @(*) begin
    pendingCmdCounter_incrementIt = 1'b0;
    if(io_input_aw_fire) begin
      pendingCmdCounter_incrementIt = 1'b1;
    end
  end

  always @(*) begin
    pendingCmdCounter_decrementIt = 1'b0;
    if(io_input_b_fire) begin
      pendingCmdCounter_decrementIt = 1'b1;
    end
  end

  assign pendingCmdCounter_willOverflowIfInc = ((pendingCmdCounter_value == 3'b111) && (! pendingCmdCounter_decrementIt));
  assign pendingCmdCounter_willOverflow = (pendingCmdCounter_willOverflowIfInc && pendingCmdCounter_incrementIt);
  assign when_Utils_l669 = (pendingCmdCounter_incrementIt && (! pendingCmdCounter_decrementIt));
  always @(*) begin
    if(when_Utils_l669) begin
      pendingCmdCounter_finalIncrement = 3'b001;
    end else begin
      if(when_Utils_l671) begin
        pendingCmdCounter_finalIncrement = 3'b111;
      end else begin
        pendingCmdCounter_finalIncrement = 3'b000;
      end
    end
  end

  assign when_Utils_l671 = ((! pendingCmdCounter_incrementIt) && pendingCmdCounter_decrementIt);
  assign pendingCmdCounter_valueNext = (pendingCmdCounter_value + pendingCmdCounter_finalIncrement);
  assign io_input_w_fire = (io_input_w_valid && io_input_w_ready);
  assign when_Utils_l644 = (io_input_w_fire && io_input_w_payload_last);
  always @(*) begin
    pendingDataCounter_incrementIt = 1'b0;
    if(cmdAllowedStart) begin
      pendingDataCounter_incrementIt = 1'b1;
    end
  end

  always @(*) begin
    pendingDataCounter_decrementIt = 1'b0;
    if(when_Utils_l644) begin
      pendingDataCounter_decrementIt = 1'b1;
    end
  end

  assign pendingDataCounter_willOverflowIfInc = ((pendingDataCounter_value == 3'b111) && (! pendingDataCounter_decrementIt));
  assign pendingDataCounter_willOverflow = (pendingDataCounter_willOverflowIfInc && pendingDataCounter_incrementIt);
  assign when_Utils_l669_1 = (pendingDataCounter_incrementIt && (! pendingDataCounter_decrementIt));
  always @(*) begin
    if(when_Utils_l669_1) begin
      pendingDataCounter_finalIncrement = 3'b001;
    end else begin
      if(when_Utils_l671_1) begin
        pendingDataCounter_finalIncrement = 3'b111;
      end else begin
        pendingDataCounter_finalIncrement = 3'b000;
      end
    end
  end

  assign when_Utils_l671_1 = ((! pendingDataCounter_incrementIt) && pendingDataCounter_decrementIt);
  assign pendingDataCounter_valueNext = (pendingDataCounter_value + pendingDataCounter_finalIncrement);
  assign decodedCmdSels = {(((32'h10000000 <= io_input_aw_payload_addr) && (io_input_aw_payload_addr < 32'h30000000)) && io_input_aw_valid),(((io_input_aw_payload_addr & (~ 32'h0001ffff)) == 32'h30000000) && io_input_aw_valid)};
  assign decodedCmdError = (decodedCmdSels == 2'b00);
  assign allowCmd = ((pendingCmdCounter_value == 3'b000) || ((pendingCmdCounter_value != 3'b111) && (pendingSels == decodedCmdSels)));
  assign allowData = (pendingDataCounter_value != 3'b000);
  assign cmdAllowedStart = ((io_input_aw_valid && allowCmd) && _zz_cmdAllowedStart);
  assign io_input_aw_ready = (((|(decodedCmdSels & {io_outputs_1_aw_ready,io_outputs_0_aw_ready})) || (decodedCmdError && errorSlave_io_axi_aw_ready)) && allowCmd);
  assign errorSlave_io_axi_aw_valid = ((io_input_aw_valid && decodedCmdError) && allowCmd);
  assign io_outputs_0_aw_valid = ((io_input_aw_valid && decodedCmdSels[0]) && allowCmd);
  assign io_outputs_0_aw_payload_addr = io_input_aw_payload_addr;
  assign io_outputs_0_aw_payload_id = io_input_aw_payload_id;
  assign io_outputs_0_aw_payload_region = io_input_aw_payload_region;
  assign io_outputs_0_aw_payload_len = io_input_aw_payload_len;
  assign io_outputs_0_aw_payload_size = io_input_aw_payload_size;
  assign io_outputs_0_aw_payload_burst = io_input_aw_payload_burst;
  assign io_outputs_0_aw_payload_lock = io_input_aw_payload_lock;
  assign io_outputs_0_aw_payload_cache = io_input_aw_payload_cache;
  assign io_outputs_0_aw_payload_qos = io_input_aw_payload_qos;
  assign io_outputs_0_aw_payload_prot = io_input_aw_payload_prot;
  assign io_outputs_1_aw_valid = ((io_input_aw_valid && decodedCmdSels[1]) && allowCmd);
  assign io_outputs_1_aw_payload_addr = io_input_aw_payload_addr;
  assign io_outputs_1_aw_payload_id = io_input_aw_payload_id;
  assign io_outputs_1_aw_payload_region = io_input_aw_payload_region;
  assign io_outputs_1_aw_payload_len = io_input_aw_payload_len;
  assign io_outputs_1_aw_payload_size = io_input_aw_payload_size;
  assign io_outputs_1_aw_payload_burst = io_input_aw_payload_burst;
  assign io_outputs_1_aw_payload_lock = io_input_aw_payload_lock;
  assign io_outputs_1_aw_payload_cache = io_input_aw_payload_cache;
  assign io_outputs_1_aw_payload_qos = io_input_aw_payload_qos;
  assign io_outputs_1_aw_payload_prot = io_input_aw_payload_prot;
  assign io_input_w_ready = (((|(pendingSels & {io_outputs_1_w_ready,io_outputs_0_w_ready})) || (pendingError && errorSlave_io_axi_w_ready)) && allowData);
  assign errorSlave_io_axi_w_valid = ((io_input_w_valid && pendingError) && allowData);
  assign _zz_io_input_b_payload_id = pendingSels[0];
  assign _zz_io_outputs_1_w_valid = pendingSels[1];
  assign io_outputs_0_w_valid = ((io_input_w_valid && _zz_io_input_b_payload_id) && allowData);
  assign io_outputs_0_w_payload_data = io_input_w_payload_data;
  assign io_outputs_0_w_payload_strb = io_input_w_payload_strb;
  assign io_outputs_0_w_payload_last = io_input_w_payload_last;
  assign io_outputs_1_w_valid = ((io_input_w_valid && _zz_io_outputs_1_w_valid) && allowData);
  assign io_outputs_1_w_payload_data = io_input_w_payload_data;
  assign io_outputs_1_w_payload_strb = io_input_w_payload_strb;
  assign io_outputs_1_w_payload_last = io_input_w_payload_last;
  assign writeRspIndex = _zz_io_outputs_1_w_valid;
  assign io_input_b_valid = ((|{io_outputs_1_b_valid,io_outputs_0_b_valid}) || errorSlave_io_axi_b_valid);
  always @(*) begin
    io_input_b_payload_id = (_zz_io_input_b_payload_id ? io_outputs_0_b_payload_id : io_outputs_1_b_payload_id);
    if(pendingError) begin
      io_input_b_payload_id = errorSlave_io_axi_b_payload_id;
    end
  end

  always @(*) begin
    io_input_b_payload_resp = (_zz_io_input_b_payload_id ? io_outputs_0_b_payload_resp : io_outputs_1_b_payload_resp);
    if(pendingError) begin
      io_input_b_payload_resp = errorSlave_io_axi_b_payload_resp;
    end
  end

  assign io_outputs_0_b_ready = io_input_b_ready;
  assign io_outputs_1_b_ready = io_input_b_ready;
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      pendingCmdCounter_value <= 3'b000;
      pendingDataCounter_value <= 3'b000;
      pendingSels <= 2'b00;
      pendingError <= 1'b0;
      _zz_cmdAllowedStart <= 1'b1;
    end else begin
      pendingCmdCounter_value <= pendingCmdCounter_valueNext;
      pendingDataCounter_value <= pendingDataCounter_valueNext;
      if(cmdAllowedStart) begin
        pendingSels <= decodedCmdSels;
      end
      if(cmdAllowedStart) begin
        pendingError <= decodedCmdError;
      end
      if(cmdAllowedStart) begin
        _zz_cmdAllowedStart <= 1'b0;
      end
      if(io_input_aw_ready) begin
        _zz_cmdAllowedStart <= 1'b1;
      end
    end
  end


endmodule

module Axi4ReadOnlyDecoder_2 (
  input               io_input_ar_valid,
  output              io_input_ar_ready,
  input      [31:0]   io_input_ar_payload_addr,
  input      [3:0]    io_input_ar_payload_id,
  input      [3:0]    io_input_ar_payload_region,
  input      [7:0]    io_input_ar_payload_len,
  input      [2:0]    io_input_ar_payload_size,
  input      [1:0]    io_input_ar_payload_burst,
  input      [0:0]    io_input_ar_payload_lock,
  input      [3:0]    io_input_ar_payload_cache,
  input      [3:0]    io_input_ar_payload_qos,
  input      [2:0]    io_input_ar_payload_prot,
  output reg          io_input_r_valid,
  input               io_input_r_ready,
  output     [31:0]   io_input_r_payload_data,
  output reg [3:0]    io_input_r_payload_id,
  output reg [1:0]    io_input_r_payload_resp,
  output reg          io_input_r_payload_last,
  output              io_outputs_0_ar_valid,
  input               io_outputs_0_ar_ready,
  output     [31:0]   io_outputs_0_ar_payload_addr,
  output     [3:0]    io_outputs_0_ar_payload_id,
  output     [3:0]    io_outputs_0_ar_payload_region,
  output     [7:0]    io_outputs_0_ar_payload_len,
  output     [2:0]    io_outputs_0_ar_payload_size,
  output     [1:0]    io_outputs_0_ar_payload_burst,
  output     [0:0]    io_outputs_0_ar_payload_lock,
  output     [3:0]    io_outputs_0_ar_payload_cache,
  output     [3:0]    io_outputs_0_ar_payload_qos,
  output     [2:0]    io_outputs_0_ar_payload_prot,
  input               io_outputs_0_r_valid,
  output              io_outputs_0_r_ready,
  input      [31:0]   io_outputs_0_r_payload_data,
  input      [3:0]    io_outputs_0_r_payload_id,
  input      [1:0]    io_outputs_0_r_payload_resp,
  input               io_outputs_0_r_payload_last,
  output              io_outputs_1_ar_valid,
  input               io_outputs_1_ar_ready,
  output     [31:0]   io_outputs_1_ar_payload_addr,
  output     [3:0]    io_outputs_1_ar_payload_id,
  output     [3:0]    io_outputs_1_ar_payload_region,
  output     [7:0]    io_outputs_1_ar_payload_len,
  output     [2:0]    io_outputs_1_ar_payload_size,
  output     [1:0]    io_outputs_1_ar_payload_burst,
  output     [0:0]    io_outputs_1_ar_payload_lock,
  output     [3:0]    io_outputs_1_ar_payload_cache,
  output     [3:0]    io_outputs_1_ar_payload_qos,
  output     [2:0]    io_outputs_1_ar_payload_prot,
  input               io_outputs_1_r_valid,
  output              io_outputs_1_r_ready,
  input      [31:0]   io_outputs_1_r_payload_data,
  input      [3:0]    io_outputs_1_r_payload_id,
  input      [1:0]    io_outputs_1_r_payload_resp,
  input               io_outputs_1_r_payload_last,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  wire                errorSlave_io_axi_ar_valid;
  wire                errorSlave_io_axi_ar_ready;
  wire                errorSlave_io_axi_r_valid;
  wire       [31:0]   errorSlave_io_axi_r_payload_data;
  wire       [3:0]    errorSlave_io_axi_r_payload_id;
  wire       [1:0]    errorSlave_io_axi_r_payload_resp;
  wire                errorSlave_io_axi_r_payload_last;
  wire                io_input_ar_fire;
  wire                io_input_r_fire;
  wire                when_Utils_l644;
  reg                 pendingCmdCounter_incrementIt;
  reg                 pendingCmdCounter_decrementIt;
  wire       [2:0]    pendingCmdCounter_valueNext;
  reg        [2:0]    pendingCmdCounter_value;
  wire                pendingCmdCounter_willOverflowIfInc;
  wire                pendingCmdCounter_willOverflow;
  reg        [2:0]    pendingCmdCounter_finalIncrement;
  wire                when_Utils_l669;
  wire                when_Utils_l671;
  wire       [1:0]    decodedCmdSels;
  wire                decodedCmdError;
  reg        [1:0]    pendingSels;
  reg                 pendingError;
  wire                allowCmd;
  wire                _zz_io_input_r_payload_data;
  wire                _zz_readRspIndex;
  wire       [0:0]    readRspIndex;

  Axi4ReadOnlyErrorSlave errorSlave (
    .io_axi_ar_valid          (errorSlave_io_axi_ar_valid            ), //i
    .io_axi_ar_ready          (errorSlave_io_axi_ar_ready            ), //o
    .io_axi_ar_payload_addr   (io_input_ar_payload_addr[31:0]        ), //i
    .io_axi_ar_payload_id     (io_input_ar_payload_id[3:0]           ), //i
    .io_axi_ar_payload_region (io_input_ar_payload_region[3:0]       ), //i
    .io_axi_ar_payload_len    (io_input_ar_payload_len[7:0]          ), //i
    .io_axi_ar_payload_size   (io_input_ar_payload_size[2:0]         ), //i
    .io_axi_ar_payload_burst  (io_input_ar_payload_burst[1:0]        ), //i
    .io_axi_ar_payload_lock   (io_input_ar_payload_lock              ), //i
    .io_axi_ar_payload_cache  (io_input_ar_payload_cache[3:0]        ), //i
    .io_axi_ar_payload_qos    (io_input_ar_payload_qos[3:0]          ), //i
    .io_axi_ar_payload_prot   (io_input_ar_payload_prot[2:0]         ), //i
    .io_axi_r_valid           (errorSlave_io_axi_r_valid             ), //o
    .io_axi_r_ready           (io_input_r_ready                      ), //i
    .io_axi_r_payload_data    (errorSlave_io_axi_r_payload_data[31:0]), //o
    .io_axi_r_payload_id      (errorSlave_io_axi_r_payload_id[3:0]   ), //o
    .io_axi_r_payload_resp    (errorSlave_io_axi_r_payload_resp[1:0] ), //o
    .io_axi_r_payload_last    (errorSlave_io_axi_r_payload_last      ), //o
    .io_axiClk                (io_axiClk                             ), //i
    .resetCtrl_axiReset       (resetCtrl_axiReset                    )  //i
  );
  assign io_input_ar_fire = (io_input_ar_valid && io_input_ar_ready);
  assign io_input_r_fire = (io_input_r_valid && io_input_r_ready);
  assign when_Utils_l644 = (io_input_r_fire && io_input_r_payload_last);
  always @(*) begin
    pendingCmdCounter_incrementIt = 1'b0;
    if(io_input_ar_fire) begin
      pendingCmdCounter_incrementIt = 1'b1;
    end
  end

  always @(*) begin
    pendingCmdCounter_decrementIt = 1'b0;
    if(when_Utils_l644) begin
      pendingCmdCounter_decrementIt = 1'b1;
    end
  end

  assign pendingCmdCounter_willOverflowIfInc = ((pendingCmdCounter_value == 3'b111) && (! pendingCmdCounter_decrementIt));
  assign pendingCmdCounter_willOverflow = (pendingCmdCounter_willOverflowIfInc && pendingCmdCounter_incrementIt);
  assign when_Utils_l669 = (pendingCmdCounter_incrementIt && (! pendingCmdCounter_decrementIt));
  always @(*) begin
    if(when_Utils_l669) begin
      pendingCmdCounter_finalIncrement = 3'b001;
    end else begin
      if(when_Utils_l671) begin
        pendingCmdCounter_finalIncrement = 3'b111;
      end else begin
        pendingCmdCounter_finalIncrement = 3'b000;
      end
    end
  end

  assign when_Utils_l671 = ((! pendingCmdCounter_incrementIt) && pendingCmdCounter_decrementIt);
  assign pendingCmdCounter_valueNext = (pendingCmdCounter_value + pendingCmdCounter_finalIncrement);
  assign decodedCmdSels = {(((32'h10000000 <= io_input_ar_payload_addr) && (io_input_ar_payload_addr < 32'h30000000)) && io_input_ar_valid),(((io_input_ar_payload_addr & (~ 32'h0001ffff)) == 32'h30000000) && io_input_ar_valid)};
  assign decodedCmdError = (decodedCmdSels == 2'b00);
  assign allowCmd = ((pendingCmdCounter_value == 3'b000) || ((pendingCmdCounter_value != 3'b111) && (pendingSels == decodedCmdSels)));
  assign io_input_ar_ready = (((|(decodedCmdSels & {io_outputs_1_ar_ready,io_outputs_0_ar_ready})) || (decodedCmdError && errorSlave_io_axi_ar_ready)) && allowCmd);
  assign errorSlave_io_axi_ar_valid = ((io_input_ar_valid && decodedCmdError) && allowCmd);
  assign io_outputs_0_ar_valid = ((io_input_ar_valid && decodedCmdSels[0]) && allowCmd);
  assign io_outputs_0_ar_payload_addr = io_input_ar_payload_addr;
  assign io_outputs_0_ar_payload_id = io_input_ar_payload_id;
  assign io_outputs_0_ar_payload_region = io_input_ar_payload_region;
  assign io_outputs_0_ar_payload_len = io_input_ar_payload_len;
  assign io_outputs_0_ar_payload_size = io_input_ar_payload_size;
  assign io_outputs_0_ar_payload_burst = io_input_ar_payload_burst;
  assign io_outputs_0_ar_payload_lock = io_input_ar_payload_lock;
  assign io_outputs_0_ar_payload_cache = io_input_ar_payload_cache;
  assign io_outputs_0_ar_payload_qos = io_input_ar_payload_qos;
  assign io_outputs_0_ar_payload_prot = io_input_ar_payload_prot;
  assign io_outputs_1_ar_valid = ((io_input_ar_valid && decodedCmdSels[1]) && allowCmd);
  assign io_outputs_1_ar_payload_addr = io_input_ar_payload_addr;
  assign io_outputs_1_ar_payload_id = io_input_ar_payload_id;
  assign io_outputs_1_ar_payload_region = io_input_ar_payload_region;
  assign io_outputs_1_ar_payload_len = io_input_ar_payload_len;
  assign io_outputs_1_ar_payload_size = io_input_ar_payload_size;
  assign io_outputs_1_ar_payload_burst = io_input_ar_payload_burst;
  assign io_outputs_1_ar_payload_lock = io_input_ar_payload_lock;
  assign io_outputs_1_ar_payload_cache = io_input_ar_payload_cache;
  assign io_outputs_1_ar_payload_qos = io_input_ar_payload_qos;
  assign io_outputs_1_ar_payload_prot = io_input_ar_payload_prot;
  assign _zz_io_input_r_payload_data = pendingSels[0];
  assign _zz_readRspIndex = pendingSels[1];
  assign readRspIndex = _zz_readRspIndex;
  always @(*) begin
    io_input_r_valid = (|{io_outputs_1_r_valid,io_outputs_0_r_valid});
    if(errorSlave_io_axi_r_valid) begin
      io_input_r_valid = 1'b1;
    end
  end

  assign io_input_r_payload_data = (_zz_io_input_r_payload_data ? io_outputs_0_r_payload_data : io_outputs_1_r_payload_data);
  always @(*) begin
    io_input_r_payload_id = (_zz_io_input_r_payload_data ? io_outputs_0_r_payload_id : io_outputs_1_r_payload_id);
    if(pendingError) begin
      io_input_r_payload_id = errorSlave_io_axi_r_payload_id;
    end
  end

  always @(*) begin
    io_input_r_payload_resp = (_zz_io_input_r_payload_data ? io_outputs_0_r_payload_resp : io_outputs_1_r_payload_resp);
    if(pendingError) begin
      io_input_r_payload_resp = errorSlave_io_axi_r_payload_resp;
    end
  end

  always @(*) begin
    io_input_r_payload_last = (_zz_io_input_r_payload_data ? io_outputs_0_r_payload_last : io_outputs_1_r_payload_last);
    if(pendingError) begin
      io_input_r_payload_last = errorSlave_io_axi_r_payload_last;
    end
  end

  assign io_outputs_0_r_ready = io_input_r_ready;
  assign io_outputs_1_r_ready = io_input_r_ready;
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      pendingCmdCounter_value <= 3'b000;
      pendingSels <= 2'b00;
      pendingError <= 1'b0;
    end else begin
      pendingCmdCounter_value <= pendingCmdCounter_valueNext;
      if(io_input_ar_ready) begin
        pendingSels <= decodedCmdSels;
      end
      if(io_input_ar_ready) begin
        pendingError <= decodedCmdError;
      end
    end
  end


endmodule

module Axi4ReadOnlyArbiter (
  input               io_inputs_0_ar_valid,
  output              io_inputs_0_ar_ready,
  input      [31:0]   io_inputs_0_ar_payload_addr,
  input      [2:0]    io_inputs_0_ar_payload_id,
  input      [3:0]    io_inputs_0_ar_payload_region,
  input      [7:0]    io_inputs_0_ar_payload_len,
  input      [2:0]    io_inputs_0_ar_payload_size,
  input      [1:0]    io_inputs_0_ar_payload_burst,
  input      [0:0]    io_inputs_0_ar_payload_lock,
  input      [3:0]    io_inputs_0_ar_payload_cache,
  input      [3:0]    io_inputs_0_ar_payload_qos,
  input      [2:0]    io_inputs_0_ar_payload_prot,
  output              io_inputs_0_r_valid,
  input               io_inputs_0_r_ready,
  output     [63:0]   io_inputs_0_r_payload_data,
  output     [2:0]    io_inputs_0_r_payload_id,
  output     [1:0]    io_inputs_0_r_payload_resp,
  output              io_inputs_0_r_payload_last,
  input               io_inputs_1_ar_valid,
  output              io_inputs_1_ar_ready,
  input      [31:0]   io_inputs_1_ar_payload_addr,
  input      [2:0]    io_inputs_1_ar_payload_id,
  input      [3:0]    io_inputs_1_ar_payload_region,
  input      [7:0]    io_inputs_1_ar_payload_len,
  input      [2:0]    io_inputs_1_ar_payload_size,
  input      [1:0]    io_inputs_1_ar_payload_burst,
  input      [0:0]    io_inputs_1_ar_payload_lock,
  input      [3:0]    io_inputs_1_ar_payload_cache,
  input      [3:0]    io_inputs_1_ar_payload_qos,
  input      [2:0]    io_inputs_1_ar_payload_prot,
  output              io_inputs_1_r_valid,
  input               io_inputs_1_r_ready,
  output     [63:0]   io_inputs_1_r_payload_data,
  output     [2:0]    io_inputs_1_r_payload_id,
  output     [1:0]    io_inputs_1_r_payload_resp,
  output              io_inputs_1_r_payload_last,
  output              io_output_ar_valid,
  input               io_output_ar_ready,
  output     [31:0]   io_output_ar_payload_addr,
  output     [3:0]    io_output_ar_payload_id,
  output     [3:0]    io_output_ar_payload_region,
  output     [7:0]    io_output_ar_payload_len,
  output     [2:0]    io_output_ar_payload_size,
  output     [1:0]    io_output_ar_payload_burst,
  output     [0:0]    io_output_ar_payload_lock,
  output     [3:0]    io_output_ar_payload_cache,
  output     [3:0]    io_output_ar_payload_qos,
  output     [2:0]    io_output_ar_payload_prot,
  input               io_output_r_valid,
  output              io_output_r_ready,
  input      [63:0]   io_output_r_payload_data,
  input      [3:0]    io_output_r_payload_id,
  input      [1:0]    io_output_r_payload_resp,
  input               io_output_r_payload_last,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  wire                cmdArbiter_io_inputs_0_ready;
  wire                cmdArbiter_io_inputs_1_ready;
  wire                cmdArbiter_io_output_valid;
  wire       [31:0]   cmdArbiter_io_output_payload_addr;
  wire       [2:0]    cmdArbiter_io_output_payload_id;
  wire       [3:0]    cmdArbiter_io_output_payload_region;
  wire       [7:0]    cmdArbiter_io_output_payload_len;
  wire       [2:0]    cmdArbiter_io_output_payload_size;
  wire       [1:0]    cmdArbiter_io_output_payload_burst;
  wire       [0:0]    cmdArbiter_io_output_payload_lock;
  wire       [3:0]    cmdArbiter_io_output_payload_cache;
  wire       [3:0]    cmdArbiter_io_output_payload_qos;
  wire       [2:0]    cmdArbiter_io_output_payload_prot;
  wire       [0:0]    cmdArbiter_io_chosen;
  wire       [1:0]    cmdArbiter_io_chosenOH;
  reg                 _zz_io_output_r_ready;
  wire       [0:0]    readRspIndex;
  wire                readRspSels_0;
  wire                readRspSels_1;

  StreamArbiter_2 cmdArbiter (
    .io_inputs_0_valid          (io_inputs_0_ar_valid                    ), //i
    .io_inputs_0_ready          (cmdArbiter_io_inputs_0_ready            ), //o
    .io_inputs_0_payload_addr   (io_inputs_0_ar_payload_addr[31:0]       ), //i
    .io_inputs_0_payload_id     (io_inputs_0_ar_payload_id[2:0]          ), //i
    .io_inputs_0_payload_region (io_inputs_0_ar_payload_region[3:0]      ), //i
    .io_inputs_0_payload_len    (io_inputs_0_ar_payload_len[7:0]         ), //i
    .io_inputs_0_payload_size   (io_inputs_0_ar_payload_size[2:0]        ), //i
    .io_inputs_0_payload_burst  (io_inputs_0_ar_payload_burst[1:0]       ), //i
    .io_inputs_0_payload_lock   (io_inputs_0_ar_payload_lock             ), //i
    .io_inputs_0_payload_cache  (io_inputs_0_ar_payload_cache[3:0]       ), //i
    .io_inputs_0_payload_qos    (io_inputs_0_ar_payload_qos[3:0]         ), //i
    .io_inputs_0_payload_prot   (io_inputs_0_ar_payload_prot[2:0]        ), //i
    .io_inputs_1_valid          (io_inputs_1_ar_valid                    ), //i
    .io_inputs_1_ready          (cmdArbiter_io_inputs_1_ready            ), //o
    .io_inputs_1_payload_addr   (io_inputs_1_ar_payload_addr[31:0]       ), //i
    .io_inputs_1_payload_id     (io_inputs_1_ar_payload_id[2:0]          ), //i
    .io_inputs_1_payload_region (io_inputs_1_ar_payload_region[3:0]      ), //i
    .io_inputs_1_payload_len    (io_inputs_1_ar_payload_len[7:0]         ), //i
    .io_inputs_1_payload_size   (io_inputs_1_ar_payload_size[2:0]        ), //i
    .io_inputs_1_payload_burst  (io_inputs_1_ar_payload_burst[1:0]       ), //i
    .io_inputs_1_payload_lock   (io_inputs_1_ar_payload_lock             ), //i
    .io_inputs_1_payload_cache  (io_inputs_1_ar_payload_cache[3:0]       ), //i
    .io_inputs_1_payload_qos    (io_inputs_1_ar_payload_qos[3:0]         ), //i
    .io_inputs_1_payload_prot   (io_inputs_1_ar_payload_prot[2:0]        ), //i
    .io_output_valid            (cmdArbiter_io_output_valid              ), //o
    .io_output_ready            (io_output_ar_ready                      ), //i
    .io_output_payload_addr     (cmdArbiter_io_output_payload_addr[31:0] ), //o
    .io_output_payload_id       (cmdArbiter_io_output_payload_id[2:0]    ), //o
    .io_output_payload_region   (cmdArbiter_io_output_payload_region[3:0]), //o
    .io_output_payload_len      (cmdArbiter_io_output_payload_len[7:0]   ), //o
    .io_output_payload_size     (cmdArbiter_io_output_payload_size[2:0]  ), //o
    .io_output_payload_burst    (cmdArbiter_io_output_payload_burst[1:0] ), //o
    .io_output_payload_lock     (cmdArbiter_io_output_payload_lock       ), //o
    .io_output_payload_cache    (cmdArbiter_io_output_payload_cache[3:0] ), //o
    .io_output_payload_qos      (cmdArbiter_io_output_payload_qos[3:0]   ), //o
    .io_output_payload_prot     (cmdArbiter_io_output_payload_prot[2:0]  ), //o
    .io_chosen                  (cmdArbiter_io_chosen                    ), //o
    .io_chosenOH                (cmdArbiter_io_chosenOH[1:0]             ), //o
    .io_axiClk                  (io_axiClk                               ), //i
    .resetCtrl_axiReset         (resetCtrl_axiReset                      )  //i
  );
  always @(*) begin
    case(readRspIndex)
      1'b0 : _zz_io_output_r_ready = io_inputs_0_r_ready;
      default : _zz_io_output_r_ready = io_inputs_1_r_ready;
    endcase
  end

  assign io_inputs_0_ar_ready = cmdArbiter_io_inputs_0_ready;
  assign io_inputs_1_ar_ready = cmdArbiter_io_inputs_1_ready;
  assign io_output_ar_valid = cmdArbiter_io_output_valid;
  assign io_output_ar_payload_addr = cmdArbiter_io_output_payload_addr;
  assign io_output_ar_payload_region = cmdArbiter_io_output_payload_region;
  assign io_output_ar_payload_len = cmdArbiter_io_output_payload_len;
  assign io_output_ar_payload_size = cmdArbiter_io_output_payload_size;
  assign io_output_ar_payload_burst = cmdArbiter_io_output_payload_burst;
  assign io_output_ar_payload_lock = cmdArbiter_io_output_payload_lock;
  assign io_output_ar_payload_cache = cmdArbiter_io_output_payload_cache;
  assign io_output_ar_payload_qos = cmdArbiter_io_output_payload_qos;
  assign io_output_ar_payload_prot = cmdArbiter_io_output_payload_prot;
  assign io_output_ar_payload_id = {cmdArbiter_io_chosen,cmdArbiter_io_output_payload_id};
  assign readRspIndex = io_output_r_payload_id[3 : 3];
  assign readRspSels_0 = (readRspIndex == 1'b0);
  assign readRspSels_1 = (readRspIndex == 1'b1);
  assign io_inputs_0_r_valid = (io_output_r_valid && readRspSels_0);
  assign io_inputs_0_r_payload_data = io_output_r_payload_data;
  assign io_inputs_0_r_payload_resp = io_output_r_payload_resp;
  assign io_inputs_0_r_payload_last = io_output_r_payload_last;
  assign io_inputs_0_r_payload_id = io_output_r_payload_id[2 : 0];
  assign io_inputs_1_r_valid = (io_output_r_valid && readRspSels_1);
  assign io_inputs_1_r_payload_data = io_output_r_payload_data;
  assign io_inputs_1_r_payload_resp = io_output_r_payload_resp;
  assign io_inputs_1_r_payload_last = io_output_r_payload_last;
  assign io_inputs_1_r_payload_id = io_output_r_payload_id[2 : 0];
  assign io_output_r_ready = _zz_io_output_r_ready;

endmodule

module Axi4SharedArbiter (
  input               io_readInputs_0_ar_valid,
  output              io_readInputs_0_ar_ready,
  input      [16:0]   io_readInputs_0_ar_payload_addr,
  input      [2:0]    io_readInputs_0_ar_payload_id,
  input      [7:0]    io_readInputs_0_ar_payload_len,
  input      [2:0]    io_readInputs_0_ar_payload_size,
  input      [1:0]    io_readInputs_0_ar_payload_burst,
  output              io_readInputs_0_r_valid,
  input               io_readInputs_0_r_ready,
  output     [63:0]   io_readInputs_0_r_payload_data,
  output     [2:0]    io_readInputs_0_r_payload_id,
  output     [1:0]    io_readInputs_0_r_payload_resp,
  output              io_readInputs_0_r_payload_last,
  input               io_readInputs_1_ar_valid,
  output              io_readInputs_1_ar_ready,
  input      [16:0]   io_readInputs_1_ar_payload_addr,
  input      [2:0]    io_readInputs_1_ar_payload_id,
  input      [7:0]    io_readInputs_1_ar_payload_len,
  input      [2:0]    io_readInputs_1_ar_payload_size,
  input      [1:0]    io_readInputs_1_ar_payload_burst,
  output              io_readInputs_1_r_valid,
  input               io_readInputs_1_r_ready,
  output     [63:0]   io_readInputs_1_r_payload_data,
  output     [2:0]    io_readInputs_1_r_payload_id,
  output     [1:0]    io_readInputs_1_r_payload_resp,
  output              io_readInputs_1_r_payload_last,
  input               io_writeInputs_0_aw_valid,
  output              io_writeInputs_0_aw_ready,
  input      [16:0]   io_writeInputs_0_aw_payload_addr,
  input      [3:0]    io_writeInputs_0_aw_payload_id,
  input      [7:0]    io_writeInputs_0_aw_payload_len,
  input      [2:0]    io_writeInputs_0_aw_payload_size,
  input      [1:0]    io_writeInputs_0_aw_payload_burst,
  input               io_writeInputs_0_w_valid,
  output              io_writeInputs_0_w_ready,
  input      [63:0]   io_writeInputs_0_w_payload_data,
  input      [7:0]    io_writeInputs_0_w_payload_strb,
  input               io_writeInputs_0_w_payload_last,
  output              io_writeInputs_0_b_valid,
  input               io_writeInputs_0_b_ready,
  output     [3:0]    io_writeInputs_0_b_payload_id,
  output     [1:0]    io_writeInputs_0_b_payload_resp,
  output              io_output_arw_valid,
  input               io_output_arw_ready,
  output     [16:0]   io_output_arw_payload_addr,
  output     [3:0]    io_output_arw_payload_id,
  output     [7:0]    io_output_arw_payload_len,
  output     [2:0]    io_output_arw_payload_size,
  output     [1:0]    io_output_arw_payload_burst,
  output              io_output_arw_payload_write,
  output              io_output_w_valid,
  input               io_output_w_ready,
  output     [63:0]   io_output_w_payload_data,
  output     [7:0]    io_output_w_payload_strb,
  output              io_output_w_payload_last,
  input               io_output_b_valid,
  output              io_output_b_ready,
  input      [3:0]    io_output_b_payload_id,
  input      [1:0]    io_output_b_payload_resp,
  input               io_output_r_valid,
  output              io_output_r_ready,
  input      [63:0]   io_output_r_payload_data,
  input      [3:0]    io_output_r_payload_id,
  input      [1:0]    io_output_r_payload_resp,
  input               io_output_r_payload_last,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  reg                 cmdArbiter_io_output_ready;
  wire                cmdRouteFork_thrown_translated_fifo_io_pop_ready;
  wire                cmdArbiter_io_inputs_0_ready;
  wire                cmdArbiter_io_inputs_1_ready;
  wire                cmdArbiter_io_inputs_2_ready;
  wire                cmdArbiter_io_output_valid;
  wire       [16:0]   cmdArbiter_io_output_payload_addr;
  wire       [2:0]    cmdArbiter_io_output_payload_id;
  wire       [7:0]    cmdArbiter_io_output_payload_len;
  wire       [2:0]    cmdArbiter_io_output_payload_size;
  wire       [1:0]    cmdArbiter_io_output_payload_burst;
  wire                cmdArbiter_io_output_payload_write;
  wire       [1:0]    cmdArbiter_io_chosen;
  wire       [2:0]    cmdArbiter_io_chosenOH;
  wire                cmdRouteFork_thrown_translated_fifo_io_push_ready;
  wire                cmdRouteFork_thrown_translated_fifo_io_pop_valid;
  wire       [2:0]    cmdRouteFork_thrown_translated_fifo_io_occupancy;
  wire       [1:0]    _zz__zz_io_output_arw_payload_id;
  wire       [3:0]    _zz_io_output_arw_payload_id_1;
  wire       [2:0]    _zz_io_output_arw_payload_id_2;
  reg                 _zz_io_output_r_ready;
  wire                inputsCmd_0_valid;
  wire                inputsCmd_0_ready;
  wire       [16:0]   inputsCmd_0_payload_addr;
  wire       [2:0]    inputsCmd_0_payload_id;
  wire       [7:0]    inputsCmd_0_payload_len;
  wire       [2:0]    inputsCmd_0_payload_size;
  wire       [1:0]    inputsCmd_0_payload_burst;
  wire                inputsCmd_0_payload_write;
  wire                inputsCmd_1_valid;
  wire                inputsCmd_1_ready;
  wire       [16:0]   inputsCmd_1_payload_addr;
  wire       [2:0]    inputsCmd_1_payload_id;
  wire       [7:0]    inputsCmd_1_payload_len;
  wire       [2:0]    inputsCmd_1_payload_size;
  wire       [1:0]    inputsCmd_1_payload_burst;
  wire                inputsCmd_1_payload_write;
  wire                inputsCmd_2_valid;
  wire                inputsCmd_2_ready;
  wire       [16:0]   inputsCmd_2_payload_addr;
  wire       [2:0]    inputsCmd_2_payload_id;
  wire       [7:0]    inputsCmd_2_payload_len;
  wire       [2:0]    inputsCmd_2_payload_size;
  wire       [1:0]    inputsCmd_2_payload_burst;
  wire                inputsCmd_2_payload_write;
  wire                cmdOutputFork_valid;
  wire                cmdOutputFork_ready;
  wire       [16:0]   cmdOutputFork_payload_addr;
  wire       [2:0]    cmdOutputFork_payload_id;
  wire       [7:0]    cmdOutputFork_payload_len;
  wire       [2:0]    cmdOutputFork_payload_size;
  wire       [1:0]    cmdOutputFork_payload_burst;
  wire                cmdOutputFork_payload_write;
  wire                cmdRouteFork_valid;
  reg                 cmdRouteFork_ready;
  wire       [16:0]   cmdRouteFork_payload_addr;
  wire       [2:0]    cmdRouteFork_payload_id;
  wire       [7:0]    cmdRouteFork_payload_len;
  wire       [2:0]    cmdRouteFork_payload_size;
  wire       [1:0]    cmdRouteFork_payload_burst;
  wire                cmdRouteFork_payload_write;
  reg                 axi_ram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_0;
  reg                 axi_ram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_1;
  wire                when_Stream_l992;
  wire                when_Stream_l992_1;
  wire                cmdOutputFork_fire;
  wire                cmdRouteFork_fire;
  wire                _zz_io_output_arw_payload_id;
  wire                when_Stream_l438;
  reg                 cmdRouteFork_thrown_valid;
  wire                cmdRouteFork_thrown_ready;
  wire       [16:0]   cmdRouteFork_thrown_payload_addr;
  wire       [2:0]    cmdRouteFork_thrown_payload_id;
  wire       [7:0]    cmdRouteFork_thrown_payload_len;
  wire       [2:0]    cmdRouteFork_thrown_payload_size;
  wire       [1:0]    cmdRouteFork_thrown_payload_burst;
  wire                cmdRouteFork_thrown_payload_write;
  wire                cmdRouteFork_thrown_translated_valid;
  wire                cmdRouteFork_thrown_translated_ready;
  wire                writeLogic_routeDataInput_valid;
  wire                writeLogic_routeDataInput_ready;
  wire       [63:0]   writeLogic_routeDataInput_payload_data;
  wire       [7:0]    writeLogic_routeDataInput_payload_strb;
  wire                writeLogic_routeDataInput_payload_last;
  wire                io_output_w_fire;
  wire                writeLogic_writeRspSels_0;
  wire       [0:0]    readRspIndex;
  wire                readRspSels_0;
  wire                readRspSels_1;

  assign _zz__zz_io_output_arw_payload_id = cmdArbiter_io_chosenOH[1 : 0];
  assign _zz_io_output_arw_payload_id_2 = cmdOutputFork_payload_id;
  assign _zz_io_output_arw_payload_id_1 = {1'd0, _zz_io_output_arw_payload_id_2};
  StreamArbiter_3 cmdArbiter (
    .io_inputs_0_valid         (inputsCmd_0_valid                      ), //i
    .io_inputs_0_ready         (cmdArbiter_io_inputs_0_ready           ), //o
    .io_inputs_0_payload_addr  (inputsCmd_0_payload_addr[16:0]         ), //i
    .io_inputs_0_payload_id    (inputsCmd_0_payload_id[2:0]            ), //i
    .io_inputs_0_payload_len   (inputsCmd_0_payload_len[7:0]           ), //i
    .io_inputs_0_payload_size  (inputsCmd_0_payload_size[2:0]          ), //i
    .io_inputs_0_payload_burst (inputsCmd_0_payload_burst[1:0]         ), //i
    .io_inputs_0_payload_write (inputsCmd_0_payload_write              ), //i
    .io_inputs_1_valid         (inputsCmd_1_valid                      ), //i
    .io_inputs_1_ready         (cmdArbiter_io_inputs_1_ready           ), //o
    .io_inputs_1_payload_addr  (inputsCmd_1_payload_addr[16:0]         ), //i
    .io_inputs_1_payload_id    (inputsCmd_1_payload_id[2:0]            ), //i
    .io_inputs_1_payload_len   (inputsCmd_1_payload_len[7:0]           ), //i
    .io_inputs_1_payload_size  (inputsCmd_1_payload_size[2:0]          ), //i
    .io_inputs_1_payload_burst (inputsCmd_1_payload_burst[1:0]         ), //i
    .io_inputs_1_payload_write (inputsCmd_1_payload_write              ), //i
    .io_inputs_2_valid         (inputsCmd_2_valid                      ), //i
    .io_inputs_2_ready         (cmdArbiter_io_inputs_2_ready           ), //o
    .io_inputs_2_payload_addr  (inputsCmd_2_payload_addr[16:0]         ), //i
    .io_inputs_2_payload_id    (inputsCmd_2_payload_id[2:0]            ), //i
    .io_inputs_2_payload_len   (inputsCmd_2_payload_len[7:0]           ), //i
    .io_inputs_2_payload_size  (inputsCmd_2_payload_size[2:0]          ), //i
    .io_inputs_2_payload_burst (inputsCmd_2_payload_burst[1:0]         ), //i
    .io_inputs_2_payload_write (inputsCmd_2_payload_write              ), //i
    .io_output_valid           (cmdArbiter_io_output_valid             ), //o
    .io_output_ready           (cmdArbiter_io_output_ready             ), //i
    .io_output_payload_addr    (cmdArbiter_io_output_payload_addr[16:0]), //o
    .io_output_payload_id      (cmdArbiter_io_output_payload_id[2:0]   ), //o
    .io_output_payload_len     (cmdArbiter_io_output_payload_len[7:0]  ), //o
    .io_output_payload_size    (cmdArbiter_io_output_payload_size[2:0] ), //o
    .io_output_payload_burst   (cmdArbiter_io_output_payload_burst[1:0]), //o
    .io_output_payload_write   (cmdArbiter_io_output_payload_write     ), //o
    .io_chosen                 (cmdArbiter_io_chosen[1:0]              ), //o
    .io_chosenOH               (cmdArbiter_io_chosenOH[2:0]            ), //o
    .io_axiClk                 (io_axiClk                              ), //i
    .resetCtrl_axiReset        (resetCtrl_axiReset                     )  //i
  );
  StreamFifoLowLatency_2 cmdRouteFork_thrown_translated_fifo (
    .io_push_valid      (cmdRouteFork_thrown_translated_valid                 ), //i
    .io_push_ready      (cmdRouteFork_thrown_translated_fifo_io_push_ready    ), //o
    .io_pop_valid       (cmdRouteFork_thrown_translated_fifo_io_pop_valid     ), //o
    .io_pop_ready       (cmdRouteFork_thrown_translated_fifo_io_pop_ready     ), //i
    .io_flush           (1'b0                                                 ), //i
    .io_occupancy       (cmdRouteFork_thrown_translated_fifo_io_occupancy[2:0]), //o
    .io_axiClk          (io_axiClk                                            ), //i
    .resetCtrl_axiReset (resetCtrl_axiReset                                   )  //i
  );
  always @(*) begin
    case(readRspIndex)
      1'b0 : _zz_io_output_r_ready = io_readInputs_0_r_ready;
      default : _zz_io_output_r_ready = io_readInputs_1_r_ready;
    endcase
  end

  assign inputsCmd_0_valid = io_readInputs_0_ar_valid;
  assign io_readInputs_0_ar_ready = inputsCmd_0_ready;
  assign inputsCmd_0_payload_addr = io_readInputs_0_ar_payload_addr;
  assign inputsCmd_0_payload_id = io_readInputs_0_ar_payload_id;
  assign inputsCmd_0_payload_len = io_readInputs_0_ar_payload_len;
  assign inputsCmd_0_payload_size = io_readInputs_0_ar_payload_size;
  assign inputsCmd_0_payload_burst = io_readInputs_0_ar_payload_burst;
  assign inputsCmd_0_payload_write = 1'b0;
  assign inputsCmd_1_valid = io_readInputs_1_ar_valid;
  assign io_readInputs_1_ar_ready = inputsCmd_1_ready;
  assign inputsCmd_1_payload_addr = io_readInputs_1_ar_payload_addr;
  assign inputsCmd_1_payload_id = io_readInputs_1_ar_payload_id;
  assign inputsCmd_1_payload_len = io_readInputs_1_ar_payload_len;
  assign inputsCmd_1_payload_size = io_readInputs_1_ar_payload_size;
  assign inputsCmd_1_payload_burst = io_readInputs_1_ar_payload_burst;
  assign inputsCmd_1_payload_write = 1'b0;
  assign inputsCmd_2_valid = io_writeInputs_0_aw_valid;
  assign io_writeInputs_0_aw_ready = inputsCmd_2_ready;
  assign inputsCmd_2_payload_addr = io_writeInputs_0_aw_payload_addr;
  assign inputsCmd_2_payload_id = io_writeInputs_0_aw_payload_id[2:0];
  assign inputsCmd_2_payload_len = io_writeInputs_0_aw_payload_len;
  assign inputsCmd_2_payload_size = io_writeInputs_0_aw_payload_size;
  assign inputsCmd_2_payload_burst = io_writeInputs_0_aw_payload_burst;
  assign inputsCmd_2_payload_write = 1'b1;
  assign inputsCmd_0_ready = cmdArbiter_io_inputs_0_ready;
  assign inputsCmd_1_ready = cmdArbiter_io_inputs_1_ready;
  assign inputsCmd_2_ready = cmdArbiter_io_inputs_2_ready;
  always @(*) begin
    cmdArbiter_io_output_ready = 1'b1;
    if(when_Stream_l992) begin
      cmdArbiter_io_output_ready = 1'b0;
    end
    if(when_Stream_l992_1) begin
      cmdArbiter_io_output_ready = 1'b0;
    end
  end

  assign when_Stream_l992 = ((! cmdOutputFork_ready) && axi_ram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_0);
  assign when_Stream_l992_1 = ((! cmdRouteFork_ready) && axi_ram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_1);
  assign cmdOutputFork_valid = (cmdArbiter_io_output_valid && axi_ram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_0);
  assign cmdOutputFork_payload_addr = cmdArbiter_io_output_payload_addr;
  assign cmdOutputFork_payload_id = cmdArbiter_io_output_payload_id;
  assign cmdOutputFork_payload_len = cmdArbiter_io_output_payload_len;
  assign cmdOutputFork_payload_size = cmdArbiter_io_output_payload_size;
  assign cmdOutputFork_payload_burst = cmdArbiter_io_output_payload_burst;
  assign cmdOutputFork_payload_write = cmdArbiter_io_output_payload_write;
  assign cmdOutputFork_fire = (cmdOutputFork_valid && cmdOutputFork_ready);
  assign cmdRouteFork_valid = (cmdArbiter_io_output_valid && axi_ram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_1);
  assign cmdRouteFork_payload_addr = cmdArbiter_io_output_payload_addr;
  assign cmdRouteFork_payload_id = cmdArbiter_io_output_payload_id;
  assign cmdRouteFork_payload_len = cmdArbiter_io_output_payload_len;
  assign cmdRouteFork_payload_size = cmdArbiter_io_output_payload_size;
  assign cmdRouteFork_payload_burst = cmdArbiter_io_output_payload_burst;
  assign cmdRouteFork_payload_write = cmdArbiter_io_output_payload_write;
  assign cmdRouteFork_fire = (cmdRouteFork_valid && cmdRouteFork_ready);
  assign io_output_arw_valid = cmdOutputFork_valid;
  assign cmdOutputFork_ready = io_output_arw_ready;
  assign io_output_arw_payload_addr = cmdOutputFork_payload_addr;
  assign io_output_arw_payload_len = cmdOutputFork_payload_len;
  assign io_output_arw_payload_size = cmdOutputFork_payload_size;
  assign io_output_arw_payload_burst = cmdOutputFork_payload_burst;
  assign io_output_arw_payload_write = cmdOutputFork_payload_write;
  assign _zz_io_output_arw_payload_id = _zz__zz_io_output_arw_payload_id[1];
  assign io_output_arw_payload_id = (cmdOutputFork_payload_write ? _zz_io_output_arw_payload_id_1 : {_zz_io_output_arw_payload_id,cmdOutputFork_payload_id});
  assign when_Stream_l438 = (! cmdRouteFork_payload_write);
  always @(*) begin
    cmdRouteFork_thrown_valid = cmdRouteFork_valid;
    if(when_Stream_l438) begin
      cmdRouteFork_thrown_valid = 1'b0;
    end
  end

  always @(*) begin
    cmdRouteFork_ready = cmdRouteFork_thrown_ready;
    if(when_Stream_l438) begin
      cmdRouteFork_ready = 1'b1;
    end
  end

  assign cmdRouteFork_thrown_payload_addr = cmdRouteFork_payload_addr;
  assign cmdRouteFork_thrown_payload_id = cmdRouteFork_payload_id;
  assign cmdRouteFork_thrown_payload_len = cmdRouteFork_payload_len;
  assign cmdRouteFork_thrown_payload_size = cmdRouteFork_payload_size;
  assign cmdRouteFork_thrown_payload_burst = cmdRouteFork_payload_burst;
  assign cmdRouteFork_thrown_payload_write = cmdRouteFork_payload_write;
  assign cmdRouteFork_thrown_translated_valid = cmdRouteFork_thrown_valid;
  assign cmdRouteFork_thrown_ready = cmdRouteFork_thrown_translated_ready;
  assign cmdRouteFork_thrown_translated_ready = cmdRouteFork_thrown_translated_fifo_io_push_ready;
  assign writeLogic_routeDataInput_valid = io_writeInputs_0_w_valid;
  assign writeLogic_routeDataInput_ready = io_writeInputs_0_w_ready;
  assign writeLogic_routeDataInput_payload_data = io_writeInputs_0_w_payload_data;
  assign writeLogic_routeDataInput_payload_strb = io_writeInputs_0_w_payload_strb;
  assign writeLogic_routeDataInput_payload_last = io_writeInputs_0_w_payload_last;
  assign io_output_w_valid = (cmdRouteFork_thrown_translated_fifo_io_pop_valid && writeLogic_routeDataInput_valid);
  assign io_output_w_payload_data = writeLogic_routeDataInput_payload_data;
  assign io_output_w_payload_strb = writeLogic_routeDataInput_payload_strb;
  assign io_output_w_payload_last = writeLogic_routeDataInput_payload_last;
  assign io_writeInputs_0_w_ready = ((cmdRouteFork_thrown_translated_fifo_io_pop_valid && io_output_w_ready) && 1'b1);
  assign io_output_w_fire = (io_output_w_valid && io_output_w_ready);
  assign cmdRouteFork_thrown_translated_fifo_io_pop_ready = (io_output_w_fire && io_output_w_payload_last);
  assign writeLogic_writeRspSels_0 = 1'b1;
  assign io_writeInputs_0_b_valid = (io_output_b_valid && writeLogic_writeRspSels_0);
  assign io_writeInputs_0_b_payload_resp = io_output_b_payload_resp;
  assign io_writeInputs_0_b_payload_id = io_output_b_payload_id;
  assign io_output_b_ready = io_writeInputs_0_b_ready;
  assign readRspIndex = io_output_r_payload_id[3 : 3];
  assign readRspSels_0 = (readRspIndex == 1'b0);
  assign readRspSels_1 = (readRspIndex == 1'b1);
  assign io_readInputs_0_r_valid = (io_output_r_valid && readRspSels_0);
  assign io_readInputs_0_r_payload_data = io_output_r_payload_data;
  assign io_readInputs_0_r_payload_resp = io_output_r_payload_resp;
  assign io_readInputs_0_r_payload_last = io_output_r_payload_last;
  assign io_readInputs_0_r_payload_id = io_output_r_payload_id[2:0];
  assign io_readInputs_1_r_valid = (io_output_r_valid && readRspSels_1);
  assign io_readInputs_1_r_payload_data = io_output_r_payload_data;
  assign io_readInputs_1_r_payload_resp = io_output_r_payload_resp;
  assign io_readInputs_1_r_payload_last = io_output_r_payload_last;
  assign io_readInputs_1_r_payload_id = io_output_r_payload_id[2:0];
  assign io_output_r_ready = _zz_io_output_r_ready;
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      axi_ram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_0 <= 1'b1;
      axi_ram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_1 <= 1'b1;
    end else begin
      if(cmdOutputFork_fire) begin
        axi_ram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_0 <= 1'b0;
      end
      if(cmdRouteFork_fire) begin
        axi_ram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_1 <= 1'b0;
      end
      if(cmdArbiter_io_output_ready) begin
        axi_ram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_0 <= 1'b1;
        axi_ram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_1 <= 1'b1;
      end
    end
  end


endmodule

module Axi4WriteOnlyDecoder (
  input               io_input_aw_valid,
  output              io_input_aw_ready,
  input      [63:0]   io_input_aw_payload_addr,
  input      [1:0]    io_input_aw_payload_id,
  input      [7:0]    io_input_aw_payload_len,
  input      [2:0]    io_input_aw_payload_size,
  input      [1:0]    io_input_aw_payload_burst,
  input               io_input_w_valid,
  output              io_input_w_ready,
  input      [63:0]   io_input_w_payload_data,
  input      [7:0]    io_input_w_payload_strb,
  input               io_input_w_payload_last,
  output              io_input_b_valid,
  input               io_input_b_ready,
  output reg [1:0]    io_input_b_payload_id,
  output reg [1:0]    io_input_b_payload_resp,
  output              io_outputs_0_aw_valid,
  input               io_outputs_0_aw_ready,
  output     [63:0]   io_outputs_0_aw_payload_addr,
  output     [1:0]    io_outputs_0_aw_payload_id,
  output     [7:0]    io_outputs_0_aw_payload_len,
  output     [2:0]    io_outputs_0_aw_payload_size,
  output     [1:0]    io_outputs_0_aw_payload_burst,
  output              io_outputs_0_w_valid,
  input               io_outputs_0_w_ready,
  output     [63:0]   io_outputs_0_w_payload_data,
  output     [7:0]    io_outputs_0_w_payload_strb,
  output              io_outputs_0_w_payload_last,
  input               io_outputs_0_b_valid,
  output              io_outputs_0_b_ready,
  input      [1:0]    io_outputs_0_b_payload_id,
  input      [1:0]    io_outputs_0_b_payload_resp,
  output              io_outputs_1_aw_valid,
  input               io_outputs_1_aw_ready,
  output     [63:0]   io_outputs_1_aw_payload_addr,
  output     [1:0]    io_outputs_1_aw_payload_id,
  output     [7:0]    io_outputs_1_aw_payload_len,
  output     [2:0]    io_outputs_1_aw_payload_size,
  output     [1:0]    io_outputs_1_aw_payload_burst,
  output              io_outputs_1_w_valid,
  input               io_outputs_1_w_ready,
  output     [63:0]   io_outputs_1_w_payload_data,
  output     [7:0]    io_outputs_1_w_payload_strb,
  output              io_outputs_1_w_payload_last,
  input               io_outputs_1_b_valid,
  output              io_outputs_1_b_ready,
  input      [1:0]    io_outputs_1_b_payload_id,
  input      [1:0]    io_outputs_1_b_payload_resp,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  wire                errorSlave_io_axi_aw_valid;
  wire                errorSlave_io_axi_w_valid;
  wire                errorSlave_io_axi_aw_ready;
  wire                errorSlave_io_axi_w_ready;
  wire                errorSlave_io_axi_b_valid;
  wire       [1:0]    errorSlave_io_axi_b_payload_id;
  wire       [1:0]    errorSlave_io_axi_b_payload_resp;
  wire                cmdAllowedStart;
  wire                io_input_aw_fire;
  wire                io_input_b_fire;
  reg                 pendingCmdCounter_incrementIt;
  reg                 pendingCmdCounter_decrementIt;
  wire       [2:0]    pendingCmdCounter_valueNext;
  reg        [2:0]    pendingCmdCounter_value;
  wire                pendingCmdCounter_willOverflowIfInc;
  wire                pendingCmdCounter_willOverflow;
  reg        [2:0]    pendingCmdCounter_finalIncrement;
  wire                when_Utils_l669;
  wire                when_Utils_l671;
  wire                io_input_w_fire;
  wire                when_Utils_l644;
  reg                 pendingDataCounter_incrementIt;
  reg                 pendingDataCounter_decrementIt;
  wire       [2:0]    pendingDataCounter_valueNext;
  reg        [2:0]    pendingDataCounter_value;
  wire                pendingDataCounter_willOverflowIfInc;
  wire                pendingDataCounter_willOverflow;
  reg        [2:0]    pendingDataCounter_finalIncrement;
  wire                when_Utils_l669_1;
  wire                when_Utils_l671_1;
  wire       [1:0]    decodedCmdSels;
  wire                decodedCmdError;
  reg        [1:0]    pendingSels;
  reg                 pendingError;
  wire                allowCmd;
  wire                allowData;
  reg                 _zz_cmdAllowedStart;
  wire                _zz_io_input_b_payload_id;
  wire                _zz_io_outputs_1_w_valid;
  wire       [0:0]    writeRspIndex;

  Axi4WriteOnlyErrorSlave_1 errorSlave (
    .io_axi_aw_valid         (errorSlave_io_axi_aw_valid           ), //i
    .io_axi_aw_ready         (errorSlave_io_axi_aw_ready           ), //o
    .io_axi_aw_payload_addr  (io_input_aw_payload_addr[63:0]       ), //i
    .io_axi_aw_payload_id    (io_input_aw_payload_id[1:0]          ), //i
    .io_axi_aw_payload_len   (io_input_aw_payload_len[7:0]         ), //i
    .io_axi_aw_payload_size  (io_input_aw_payload_size[2:0]        ), //i
    .io_axi_aw_payload_burst (io_input_aw_payload_burst[1:0]       ), //i
    .io_axi_w_valid          (errorSlave_io_axi_w_valid            ), //i
    .io_axi_w_ready          (errorSlave_io_axi_w_ready            ), //o
    .io_axi_w_payload_data   (io_input_w_payload_data[63:0]        ), //i
    .io_axi_w_payload_strb   (io_input_w_payload_strb[7:0]         ), //i
    .io_axi_w_payload_last   (io_input_w_payload_last              ), //i
    .io_axi_b_valid          (errorSlave_io_axi_b_valid            ), //o
    .io_axi_b_ready          (io_input_b_ready                     ), //i
    .io_axi_b_payload_id     (errorSlave_io_axi_b_payload_id[1:0]  ), //o
    .io_axi_b_payload_resp   (errorSlave_io_axi_b_payload_resp[1:0]), //o
    .io_axiClk               (io_axiClk                            ), //i
    .resetCtrl_axiReset      (resetCtrl_axiReset                   )  //i
  );
  assign io_input_aw_fire = (io_input_aw_valid && io_input_aw_ready);
  assign io_input_b_fire = (io_input_b_valid && io_input_b_ready);
  always @(*) begin
    pendingCmdCounter_incrementIt = 1'b0;
    if(io_input_aw_fire) begin
      pendingCmdCounter_incrementIt = 1'b1;
    end
  end

  always @(*) begin
    pendingCmdCounter_decrementIt = 1'b0;
    if(io_input_b_fire) begin
      pendingCmdCounter_decrementIt = 1'b1;
    end
  end

  assign pendingCmdCounter_willOverflowIfInc = ((pendingCmdCounter_value == 3'b111) && (! pendingCmdCounter_decrementIt));
  assign pendingCmdCounter_willOverflow = (pendingCmdCounter_willOverflowIfInc && pendingCmdCounter_incrementIt);
  assign when_Utils_l669 = (pendingCmdCounter_incrementIt && (! pendingCmdCounter_decrementIt));
  always @(*) begin
    if(when_Utils_l669) begin
      pendingCmdCounter_finalIncrement = 3'b001;
    end else begin
      if(when_Utils_l671) begin
        pendingCmdCounter_finalIncrement = 3'b111;
      end else begin
        pendingCmdCounter_finalIncrement = 3'b000;
      end
    end
  end

  assign when_Utils_l671 = ((! pendingCmdCounter_incrementIt) && pendingCmdCounter_decrementIt);
  assign pendingCmdCounter_valueNext = (pendingCmdCounter_value + pendingCmdCounter_finalIncrement);
  assign io_input_w_fire = (io_input_w_valid && io_input_w_ready);
  assign when_Utils_l644 = (io_input_w_fire && io_input_w_payload_last);
  always @(*) begin
    pendingDataCounter_incrementIt = 1'b0;
    if(cmdAllowedStart) begin
      pendingDataCounter_incrementIt = 1'b1;
    end
  end

  always @(*) begin
    pendingDataCounter_decrementIt = 1'b0;
    if(when_Utils_l644) begin
      pendingDataCounter_decrementIt = 1'b1;
    end
  end

  assign pendingDataCounter_willOverflowIfInc = ((pendingDataCounter_value == 3'b111) && (! pendingDataCounter_decrementIt));
  assign pendingDataCounter_willOverflow = (pendingDataCounter_willOverflowIfInc && pendingDataCounter_incrementIt);
  assign when_Utils_l669_1 = (pendingDataCounter_incrementIt && (! pendingDataCounter_decrementIt));
  always @(*) begin
    if(when_Utils_l669_1) begin
      pendingDataCounter_finalIncrement = 3'b001;
    end else begin
      if(when_Utils_l671_1) begin
        pendingDataCounter_finalIncrement = 3'b111;
      end else begin
        pendingDataCounter_finalIncrement = 3'b000;
      end
    end
  end

  assign when_Utils_l671_1 = ((! pendingDataCounter_incrementIt) && pendingDataCounter_decrementIt);
  assign pendingDataCounter_valueNext = (pendingDataCounter_value + pendingDataCounter_finalIncrement);
  assign decodedCmdSels = {(((64'h0000000010000000 <= io_input_aw_payload_addr) && (io_input_aw_payload_addr < 64'h0000000040000000)) && io_input_aw_valid),(((io_input_aw_payload_addr & (~ 64'h000000000001ffff)) == 64'h0000000080000000) && io_input_aw_valid)};
  assign decodedCmdError = (decodedCmdSels == 2'b00);
  assign allowCmd = ((pendingCmdCounter_value == 3'b000) || ((pendingCmdCounter_value != 3'b111) && (pendingSels == decodedCmdSels)));
  assign allowData = (pendingDataCounter_value != 3'b000);
  assign cmdAllowedStart = ((io_input_aw_valid && allowCmd) && _zz_cmdAllowedStart);
  assign io_input_aw_ready = (((|(decodedCmdSels & {io_outputs_1_aw_ready,io_outputs_0_aw_ready})) || (decodedCmdError && errorSlave_io_axi_aw_ready)) && allowCmd);
  assign errorSlave_io_axi_aw_valid = ((io_input_aw_valid && decodedCmdError) && allowCmd);
  assign io_outputs_0_aw_valid = ((io_input_aw_valid && decodedCmdSels[0]) && allowCmd);
  assign io_outputs_0_aw_payload_addr = io_input_aw_payload_addr;
  assign io_outputs_0_aw_payload_id = io_input_aw_payload_id;
  assign io_outputs_0_aw_payload_len = io_input_aw_payload_len;
  assign io_outputs_0_aw_payload_size = io_input_aw_payload_size;
  assign io_outputs_0_aw_payload_burst = io_input_aw_payload_burst;
  assign io_outputs_1_aw_valid = ((io_input_aw_valid && decodedCmdSels[1]) && allowCmd);
  assign io_outputs_1_aw_payload_addr = io_input_aw_payload_addr;
  assign io_outputs_1_aw_payload_id = io_input_aw_payload_id;
  assign io_outputs_1_aw_payload_len = io_input_aw_payload_len;
  assign io_outputs_1_aw_payload_size = io_input_aw_payload_size;
  assign io_outputs_1_aw_payload_burst = io_input_aw_payload_burst;
  assign io_input_w_ready = (((|(pendingSels & {io_outputs_1_w_ready,io_outputs_0_w_ready})) || (pendingError && errorSlave_io_axi_w_ready)) && allowData);
  assign errorSlave_io_axi_w_valid = ((io_input_w_valid && pendingError) && allowData);
  assign _zz_io_input_b_payload_id = pendingSels[0];
  assign _zz_io_outputs_1_w_valid = pendingSels[1];
  assign io_outputs_0_w_valid = ((io_input_w_valid && _zz_io_input_b_payload_id) && allowData);
  assign io_outputs_0_w_payload_data = io_input_w_payload_data;
  assign io_outputs_0_w_payload_strb = io_input_w_payload_strb;
  assign io_outputs_0_w_payload_last = io_input_w_payload_last;
  assign io_outputs_1_w_valid = ((io_input_w_valid && _zz_io_outputs_1_w_valid) && allowData);
  assign io_outputs_1_w_payload_data = io_input_w_payload_data;
  assign io_outputs_1_w_payload_strb = io_input_w_payload_strb;
  assign io_outputs_1_w_payload_last = io_input_w_payload_last;
  assign writeRspIndex = _zz_io_outputs_1_w_valid;
  assign io_input_b_valid = ((|{io_outputs_1_b_valid,io_outputs_0_b_valid}) || errorSlave_io_axi_b_valid);
  always @(*) begin
    io_input_b_payload_id = (_zz_io_input_b_payload_id ? io_outputs_0_b_payload_id : io_outputs_1_b_payload_id);
    if(pendingError) begin
      io_input_b_payload_id = errorSlave_io_axi_b_payload_id;
    end
  end

  always @(*) begin
    io_input_b_payload_resp = (_zz_io_input_b_payload_id ? io_outputs_0_b_payload_resp : io_outputs_1_b_payload_resp);
    if(pendingError) begin
      io_input_b_payload_resp = errorSlave_io_axi_b_payload_resp;
    end
  end

  assign io_outputs_0_b_ready = io_input_b_ready;
  assign io_outputs_1_b_ready = io_input_b_ready;
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      pendingCmdCounter_value <= 3'b000;
      pendingDataCounter_value <= 3'b000;
      pendingSels <= 2'b00;
      pendingError <= 1'b0;
      _zz_cmdAllowedStart <= 1'b1;
    end else begin
      pendingCmdCounter_value <= pendingCmdCounter_valueNext;
      pendingDataCounter_value <= pendingDataCounter_valueNext;
      if(cmdAllowedStart) begin
        pendingSels <= decodedCmdSels;
      end
      if(cmdAllowedStart) begin
        pendingError <= decodedCmdError;
      end
      if(cmdAllowedStart) begin
        _zz_cmdAllowedStart <= 1'b0;
      end
      if(io_input_aw_ready) begin
        _zz_cmdAllowedStart <= 1'b1;
      end
    end
  end


endmodule

//Axi4ReadOnlyDecoder_1 replaced by Axi4ReadOnlyDecoder

module Axi4ReadOnlyDecoder (
  input               io_input_ar_valid,
  output              io_input_ar_ready,
  input      [63:0]   io_input_ar_payload_addr,
  input      [1:0]    io_input_ar_payload_id,
  input      [7:0]    io_input_ar_payload_len,
  input      [2:0]    io_input_ar_payload_size,
  input      [1:0]    io_input_ar_payload_burst,
  output reg          io_input_r_valid,
  input               io_input_r_ready,
  output     [63:0]   io_input_r_payload_data,
  output reg [1:0]    io_input_r_payload_id,
  output reg [1:0]    io_input_r_payload_resp,
  output reg          io_input_r_payload_last,
  output              io_outputs_0_ar_valid,
  input               io_outputs_0_ar_ready,
  output     [63:0]   io_outputs_0_ar_payload_addr,
  output     [1:0]    io_outputs_0_ar_payload_id,
  output     [7:0]    io_outputs_0_ar_payload_len,
  output     [2:0]    io_outputs_0_ar_payload_size,
  output     [1:0]    io_outputs_0_ar_payload_burst,
  input               io_outputs_0_r_valid,
  output              io_outputs_0_r_ready,
  input      [63:0]   io_outputs_0_r_payload_data,
  input      [1:0]    io_outputs_0_r_payload_id,
  input      [1:0]    io_outputs_0_r_payload_resp,
  input               io_outputs_0_r_payload_last,
  output              io_outputs_1_ar_valid,
  input               io_outputs_1_ar_ready,
  output     [63:0]   io_outputs_1_ar_payload_addr,
  output     [1:0]    io_outputs_1_ar_payload_id,
  output     [7:0]    io_outputs_1_ar_payload_len,
  output     [2:0]    io_outputs_1_ar_payload_size,
  output     [1:0]    io_outputs_1_ar_payload_burst,
  input               io_outputs_1_r_valid,
  output              io_outputs_1_r_ready,
  input      [63:0]   io_outputs_1_r_payload_data,
  input      [1:0]    io_outputs_1_r_payload_id,
  input      [1:0]    io_outputs_1_r_payload_resp,
  input               io_outputs_1_r_payload_last,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  wire                errorSlave_io_axi_ar_valid;
  wire                errorSlave_io_axi_ar_ready;
  wire                errorSlave_io_axi_r_valid;
  wire       [63:0]   errorSlave_io_axi_r_payload_data;
  wire       [1:0]    errorSlave_io_axi_r_payload_id;
  wire       [1:0]    errorSlave_io_axi_r_payload_resp;
  wire                errorSlave_io_axi_r_payload_last;
  wire                io_input_ar_fire;
  wire                io_input_r_fire;
  wire                when_Utils_l644;
  reg                 pendingCmdCounter_incrementIt;
  reg                 pendingCmdCounter_decrementIt;
  wire       [2:0]    pendingCmdCounter_valueNext;
  reg        [2:0]    pendingCmdCounter_value;
  wire                pendingCmdCounter_willOverflowIfInc;
  wire                pendingCmdCounter_willOverflow;
  reg        [2:0]    pendingCmdCounter_finalIncrement;
  wire                when_Utils_l669;
  wire                when_Utils_l671;
  wire       [1:0]    decodedCmdSels;
  wire                decodedCmdError;
  reg        [1:0]    pendingSels;
  reg                 pendingError;
  wire                allowCmd;
  wire                _zz_io_input_r_payload_data;
  wire                _zz_readRspIndex;
  wire       [0:0]    readRspIndex;

  Axi4ReadOnlyErrorSlave_2 errorSlave (
    .io_axi_ar_valid         (errorSlave_io_axi_ar_valid            ), //i
    .io_axi_ar_ready         (errorSlave_io_axi_ar_ready            ), //o
    .io_axi_ar_payload_addr  (io_input_ar_payload_addr[63:0]        ), //i
    .io_axi_ar_payload_id    (io_input_ar_payload_id[1:0]           ), //i
    .io_axi_ar_payload_len   (io_input_ar_payload_len[7:0]          ), //i
    .io_axi_ar_payload_size  (io_input_ar_payload_size[2:0]         ), //i
    .io_axi_ar_payload_burst (io_input_ar_payload_burst[1:0]        ), //i
    .io_axi_r_valid          (errorSlave_io_axi_r_valid             ), //o
    .io_axi_r_ready          (io_input_r_ready                      ), //i
    .io_axi_r_payload_data   (errorSlave_io_axi_r_payload_data[63:0]), //o
    .io_axi_r_payload_id     (errorSlave_io_axi_r_payload_id[1:0]   ), //o
    .io_axi_r_payload_resp   (errorSlave_io_axi_r_payload_resp[1:0] ), //o
    .io_axi_r_payload_last   (errorSlave_io_axi_r_payload_last      ), //o
    .io_axiClk               (io_axiClk                             ), //i
    .resetCtrl_axiReset      (resetCtrl_axiReset                    )  //i
  );
  assign io_input_ar_fire = (io_input_ar_valid && io_input_ar_ready);
  assign io_input_r_fire = (io_input_r_valid && io_input_r_ready);
  assign when_Utils_l644 = (io_input_r_fire && io_input_r_payload_last);
  always @(*) begin
    pendingCmdCounter_incrementIt = 1'b0;
    if(io_input_ar_fire) begin
      pendingCmdCounter_incrementIt = 1'b1;
    end
  end

  always @(*) begin
    pendingCmdCounter_decrementIt = 1'b0;
    if(when_Utils_l644) begin
      pendingCmdCounter_decrementIt = 1'b1;
    end
  end

  assign pendingCmdCounter_willOverflowIfInc = ((pendingCmdCounter_value == 3'b111) && (! pendingCmdCounter_decrementIt));
  assign pendingCmdCounter_willOverflow = (pendingCmdCounter_willOverflowIfInc && pendingCmdCounter_incrementIt);
  assign when_Utils_l669 = (pendingCmdCounter_incrementIt && (! pendingCmdCounter_decrementIt));
  always @(*) begin
    if(when_Utils_l669) begin
      pendingCmdCounter_finalIncrement = 3'b001;
    end else begin
      if(when_Utils_l671) begin
        pendingCmdCounter_finalIncrement = 3'b111;
      end else begin
        pendingCmdCounter_finalIncrement = 3'b000;
      end
    end
  end

  assign when_Utils_l671 = ((! pendingCmdCounter_incrementIt) && pendingCmdCounter_decrementIt);
  assign pendingCmdCounter_valueNext = (pendingCmdCounter_value + pendingCmdCounter_finalIncrement);
  assign decodedCmdSels = {(((64'h0000000010000000 <= io_input_ar_payload_addr) && (io_input_ar_payload_addr < 64'h0000000040000000)) && io_input_ar_valid),(((io_input_ar_payload_addr & (~ 64'h000000000001ffff)) == 64'h0000000080000000) && io_input_ar_valid)};
  assign decodedCmdError = (decodedCmdSels == 2'b00);
  assign allowCmd = ((pendingCmdCounter_value == 3'b000) || ((pendingCmdCounter_value != 3'b111) && (pendingSels == decodedCmdSels)));
  assign io_input_ar_ready = (((|(decodedCmdSels & {io_outputs_1_ar_ready,io_outputs_0_ar_ready})) || (decodedCmdError && errorSlave_io_axi_ar_ready)) && allowCmd);
  assign errorSlave_io_axi_ar_valid = ((io_input_ar_valid && decodedCmdError) && allowCmd);
  assign io_outputs_0_ar_valid = ((io_input_ar_valid && decodedCmdSels[0]) && allowCmd);
  assign io_outputs_0_ar_payload_addr = io_input_ar_payload_addr;
  assign io_outputs_0_ar_payload_id = io_input_ar_payload_id;
  assign io_outputs_0_ar_payload_len = io_input_ar_payload_len;
  assign io_outputs_0_ar_payload_size = io_input_ar_payload_size;
  assign io_outputs_0_ar_payload_burst = io_input_ar_payload_burst;
  assign io_outputs_1_ar_valid = ((io_input_ar_valid && decodedCmdSels[1]) && allowCmd);
  assign io_outputs_1_ar_payload_addr = io_input_ar_payload_addr;
  assign io_outputs_1_ar_payload_id = io_input_ar_payload_id;
  assign io_outputs_1_ar_payload_len = io_input_ar_payload_len;
  assign io_outputs_1_ar_payload_size = io_input_ar_payload_size;
  assign io_outputs_1_ar_payload_burst = io_input_ar_payload_burst;
  assign _zz_io_input_r_payload_data = pendingSels[0];
  assign _zz_readRspIndex = pendingSels[1];
  assign readRspIndex = _zz_readRspIndex;
  always @(*) begin
    io_input_r_valid = (|{io_outputs_1_r_valid,io_outputs_0_r_valid});
    if(errorSlave_io_axi_r_valid) begin
      io_input_r_valid = 1'b1;
    end
  end

  assign io_input_r_payload_data = (_zz_io_input_r_payload_data ? io_outputs_0_r_payload_data : io_outputs_1_r_payload_data);
  always @(*) begin
    io_input_r_payload_id = (_zz_io_input_r_payload_data ? io_outputs_0_r_payload_id : io_outputs_1_r_payload_id);
    if(pendingError) begin
      io_input_r_payload_id = errorSlave_io_axi_r_payload_id;
    end
  end

  always @(*) begin
    io_input_r_payload_resp = (_zz_io_input_r_payload_data ? io_outputs_0_r_payload_resp : io_outputs_1_r_payload_resp);
    if(pendingError) begin
      io_input_r_payload_resp = errorSlave_io_axi_r_payload_resp;
    end
  end

  always @(*) begin
    io_input_r_payload_last = (_zz_io_input_r_payload_data ? io_outputs_0_r_payload_last : io_outputs_1_r_payload_last);
    if(pendingError) begin
      io_input_r_payload_last = errorSlave_io_axi_r_payload_last;
    end
  end

  assign io_outputs_0_r_ready = io_input_r_ready;
  assign io_outputs_1_r_ready = io_input_r_ready;
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      pendingCmdCounter_value <= 3'b000;
      pendingSels <= 2'b00;
      pendingError <= 1'b0;
    end else begin
      pendingCmdCounter_value <= pendingCmdCounter_valueNext;
      if(io_input_ar_ready) begin
        pendingSels <= decodedCmdSels;
      end
      if(io_input_ar_ready) begin
        pendingError <= decodedCmdError;
      end
    end
  end


endmodule

module Apb3Uart (
  input      [15:0]   io_apb_PADDR /* verilator public */ ,
  input      [0:0]    io_apb_PSEL /* verilator public */ ,
  input               io_apb_PENABLE /* verilator public */ ,
  output              io_apb_PREADY /* verilator public */ ,
  input               io_apb_PWRITE /* verilator public */ ,
  input      [31:0]   io_apb_PWDATA /* verilator public */ ,
  output     [31:0]   io_apb_PRDATA /* verilator public */ ,
  output              io_apb_PSLVERROR /* verilator public */ ,
  output              io_uart_txd,
  input               io_uart_rxd,
  input               io_clock,
  input               io_resetn
);

  wire       [31:0]   uartCtrl_in_paddr;
  wire                uartCtrl_in_pwrite;
  wire                uartCtrl_in_pready;
  wire                uartCtrl_in_pslverr;
  wire       [31:0]   uartCtrl_in_prdata;
  wire                uartCtrl_uart_tx;

  uart_apb uartCtrl (
    .clk        (io_clock                ), //i
    .resetn     (io_resetn               ), //i
    .in_psel    (io_apb_PSEL             ), //i
    .in_penable (io_apb_PENABLE          ), //i
    .in_pprot   (3'b000                  ), //i
    .in_pready  (uartCtrl_in_pready      ), //o
    .in_pslverr (uartCtrl_in_pslverr     ), //o
    .in_paddr   (uartCtrl_in_paddr[31:0] ), //i
    .in_pwrite  (uartCtrl_in_pwrite      ), //i
    .in_prdata  (uartCtrl_in_prdata[31:0]), //o
    .in_pwdata  (io_apb_PWDATA[31:0]     ), //i
    .in_pstrb   (4'b1111                 ), //i
    .uart_rx    (io_uart_rxd             ), //i
    .uart_tx    (uartCtrl_uart_tx        )  //o
  );
  assign io_uart_txd = uartCtrl_uart_tx;
  assign io_apb_PREADY = uartCtrl_in_pready;
  assign io_apb_PSLVERROR = uartCtrl_in_pslverr;
  assign uartCtrl_in_paddr = {16'd0, io_apb_PADDR};
  assign uartCtrl_in_pwrite = ((io_apb_PWRITE && io_apb_PENABLE) && io_apb_PSEL[0]);
  assign io_apb_PRDATA = uartCtrl_in_prdata;

endmodule

module Axi4SharedToApb3Bridge (
  input               io_axi_arw_valid,
  output reg          io_axi_arw_ready,
  input      [19:0]   io_axi_arw_payload_addr,
  input      [3:0]    io_axi_arw_payload_id,
  input      [7:0]    io_axi_arw_payload_len,
  input      [2:0]    io_axi_arw_payload_size,
  input      [1:0]    io_axi_arw_payload_burst,
  input               io_axi_arw_payload_write,
  input               io_axi_w_valid,
  output reg          io_axi_w_ready,
  input      [31:0]   io_axi_w_payload_data,
  input      [3:0]    io_axi_w_payload_strb,
  input               io_axi_w_payload_last,
  output reg          io_axi_b_valid,
  input               io_axi_b_ready,
  output     [3:0]    io_axi_b_payload_id,
  output     [1:0]    io_axi_b_payload_resp,
  output reg          io_axi_r_valid,
  input               io_axi_r_ready,
  output     [31:0]   io_axi_r_payload_data,
  output     [3:0]    io_axi_r_payload_id,
  output     [1:0]    io_axi_r_payload_resp,
  output              io_axi_r_payload_last,
  output     [19:0]   io_apb_PADDR,
  output reg [0:0]    io_apb_PSEL,
  output reg          io_apb_PENABLE,
  input               io_apb_PREADY,
  output              io_apb_PWRITE,
  output     [31:0]   io_apb_PWDATA,
  input      [31:0]   io_apb_PRDATA,
  input               io_apb_PSLVERROR,
  input               io_axiClk,
  input               resetCtrl_axiReset
);
  localparam Axi4ToApb3BridgePhase_SETUP = 2'd0;
  localparam Axi4ToApb3BridgePhase_ACCESS_1 = 2'd1;
  localparam Axi4ToApb3BridgePhase_RESPONSE = 2'd2;

  reg        [1:0]    phase;
  reg                 write;
  reg        [31:0]   readedData;
  reg        [3:0]    id;
  wire                when_Axi4SharedToApb3Bridge_l91;
  wire                when_Axi4SharedToApb3Bridge_l97;
  `ifndef SYNTHESIS
  reg [63:0] phase_string;
  `endif


  `ifndef SYNTHESIS
  always @(*) begin
    case(phase)
      Axi4ToApb3BridgePhase_SETUP : phase_string = "SETUP   ";
      Axi4ToApb3BridgePhase_ACCESS_1 : phase_string = "ACCESS_1";
      Axi4ToApb3BridgePhase_RESPONSE : phase_string = "RESPONSE";
      default : phase_string = "????????";
    endcase
  end
  `endif

  always @(*) begin
    io_axi_arw_ready = 1'b0;
    case(phase)
      Axi4ToApb3BridgePhase_SETUP : begin
        if(when_Axi4SharedToApb3Bridge_l91) begin
          if(when_Axi4SharedToApb3Bridge_l97) begin
            io_axi_arw_ready = 1'b1;
          end
        end
      end
      Axi4ToApb3BridgePhase_ACCESS_1 : begin
        if(io_apb_PREADY) begin
          io_axi_arw_ready = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axi_w_ready = 1'b0;
    case(phase)
      Axi4ToApb3BridgePhase_SETUP : begin
        if(when_Axi4SharedToApb3Bridge_l91) begin
          if(when_Axi4SharedToApb3Bridge_l97) begin
            io_axi_w_ready = 1'b1;
          end
        end
      end
      Axi4ToApb3BridgePhase_ACCESS_1 : begin
        if(io_apb_PREADY) begin
          io_axi_w_ready = write;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axi_b_valid = 1'b0;
    case(phase)
      Axi4ToApb3BridgePhase_SETUP : begin
      end
      Axi4ToApb3BridgePhase_ACCESS_1 : begin
      end
      default : begin
        if(write) begin
          io_axi_b_valid = 1'b1;
        end
      end
    endcase
  end

  always @(*) begin
    io_axi_r_valid = 1'b0;
    case(phase)
      Axi4ToApb3BridgePhase_SETUP : begin
      end
      Axi4ToApb3BridgePhase_ACCESS_1 : begin
      end
      default : begin
        if(!write) begin
          io_axi_r_valid = 1'b1;
        end
      end
    endcase
  end

  always @(*) begin
    io_apb_PSEL[0] = 1'b0;
    case(phase)
      Axi4ToApb3BridgePhase_SETUP : begin
        if(when_Axi4SharedToApb3Bridge_l91) begin
          io_apb_PSEL[0] = 1'b1;
          if(when_Axi4SharedToApb3Bridge_l97) begin
            io_apb_PSEL[0] = 1'b0;
          end
        end
      end
      Axi4ToApb3BridgePhase_ACCESS_1 : begin
        io_apb_PSEL[0] = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_apb_PENABLE = 1'b0;
    case(phase)
      Axi4ToApb3BridgePhase_SETUP : begin
      end
      Axi4ToApb3BridgePhase_ACCESS_1 : begin
        io_apb_PENABLE = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign when_Axi4SharedToApb3Bridge_l91 = (io_axi_arw_valid && ((! io_axi_arw_payload_write) || io_axi_w_valid));
  assign when_Axi4SharedToApb3Bridge_l97 = (io_axi_arw_payload_write && (io_axi_w_payload_strb == 4'b0000));
  assign io_apb_PADDR = io_axi_arw_payload_addr;
  assign io_apb_PWDATA = io_axi_w_payload_data;
  assign io_apb_PWRITE = io_axi_arw_payload_write;
  assign io_axi_r_payload_resp = {io_apb_PSLVERROR,1'b0};
  assign io_axi_b_payload_resp = {io_apb_PSLVERROR,1'b0};
  assign io_axi_r_payload_id = id;
  assign io_axi_b_payload_id = id;
  assign io_axi_r_payload_data = readedData;
  assign io_axi_r_payload_last = 1'b1;
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      phase <= Axi4ToApb3BridgePhase_SETUP;
    end else begin
      case(phase)
        Axi4ToApb3BridgePhase_SETUP : begin
          if(when_Axi4SharedToApb3Bridge_l91) begin
            phase <= Axi4ToApb3BridgePhase_ACCESS_1;
            if(when_Axi4SharedToApb3Bridge_l97) begin
              phase <= Axi4ToApb3BridgePhase_RESPONSE;
            end
          end
        end
        Axi4ToApb3BridgePhase_ACCESS_1 : begin
          if(io_apb_PREADY) begin
            phase <= Axi4ToApb3BridgePhase_RESPONSE;
          end
        end
        default : begin
          if(write) begin
            if(io_axi_b_ready) begin
              phase <= Axi4ToApb3BridgePhase_SETUP;
            end
          end else begin
            if(io_axi_r_ready) begin
              phase <= Axi4ToApb3BridgePhase_SETUP;
            end
          end
        end
      endcase
    end
  end

  always @(posedge io_axiClk) begin
    case(phase)
      Axi4ToApb3BridgePhase_SETUP : begin
        write <= io_axi_arw_payload_write;
        id <= io_axi_arw_payload_id;
      end
      Axi4ToApb3BridgePhase_ACCESS_1 : begin
        if(io_apb_PREADY) begin
          readedData <= io_apb_PRDATA;
        end
      end
      default : begin
      end
    endcase
  end


endmodule

module Axi4SharedOnChipRam_1 (
  input               io_axi_arw_valid,
  output reg          io_axi_arw_ready,
  input      [16:0]   io_axi_arw_payload_addr,
  input      [3:0]    io_axi_arw_payload_id,
  input      [7:0]    io_axi_arw_payload_len,
  input      [2:0]    io_axi_arw_payload_size,
  input      [1:0]    io_axi_arw_payload_burst,
  input               io_axi_arw_payload_write,
  input               io_axi_w_valid,
  output              io_axi_w_ready,
  input      [31:0]   io_axi_w_payload_data,
  input      [3:0]    io_axi_w_payload_strb,
  input               io_axi_w_payload_last,
  output              io_axi_b_valid,
  input               io_axi_b_ready,
  output     [3:0]    io_axi_b_payload_id,
  output     [1:0]    io_axi_b_payload_resp,
  output              io_axi_r_valid,
  input               io_axi_r_ready,
  output     [31:0]   io_axi_r_payload_data,
  output     [3:0]    io_axi_r_payload_id,
  output     [1:0]    io_axi_r_payload_resp,
  output              io_axi_r_payload_last,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  reg        [31:0]   _zz_ram_port0;
  wire       [1:0]    _zz_Axi4Incr_alignMask;
  wire       [11:0]   _zz_Axi4Incr_base;
  wire       [11:0]   _zz_Axi4Incr_base_1;
  wire       [11:0]   _zz_Axi4Incr_baseIncr;
  wire       [2:0]    _zz_Axi4Incr_wrapCase_1;
  wire       [2:0]    _zz_Axi4Incr_wrapCase_2;
  reg        [11:0]   _zz_Axi4Incr_result;
  wire       [10:0]   _zz_Axi4Incr_result_1;
  wire       [0:0]    _zz_Axi4Incr_result_2;
  wire       [9:0]    _zz_Axi4Incr_result_3;
  wire       [1:0]    _zz_Axi4Incr_result_4;
  wire       [8:0]    _zz_Axi4Incr_result_5;
  wire       [2:0]    _zz_Axi4Incr_result_6;
  wire       [7:0]    _zz_Axi4Incr_result_7;
  wire       [3:0]    _zz_Axi4Incr_result_8;
  wire       [6:0]    _zz_Axi4Incr_result_9;
  wire       [4:0]    _zz_Axi4Incr_result_10;
  wire       [5:0]    _zz_Axi4Incr_result_11;
  wire       [5:0]    _zz_Axi4Incr_result_12;
  reg                 unburstify_result_valid;
  wire                unburstify_result_ready;
  reg                 unburstify_result_payload_last;
  reg        [16:0]   unburstify_result_payload_fragment_addr;
  reg        [3:0]    unburstify_result_payload_fragment_id;
  reg        [2:0]    unburstify_result_payload_fragment_size;
  reg        [1:0]    unburstify_result_payload_fragment_burst;
  reg                 unburstify_result_payload_fragment_write;
  wire                unburstify_doResult;
  reg                 unburstify_buffer_valid;
  reg        [7:0]    unburstify_buffer_len;
  reg        [7:0]    unburstify_buffer_beat;
  reg        [16:0]   unburstify_buffer_transaction_addr;
  reg        [3:0]    unburstify_buffer_transaction_id;
  reg        [2:0]    unburstify_buffer_transaction_size;
  reg        [1:0]    unburstify_buffer_transaction_burst;
  reg                 unburstify_buffer_transaction_write;
  wire                unburstify_buffer_last;
  wire       [1:0]    Axi4Incr_validSize;
  reg        [16:0]   Axi4Incr_result;
  wire       [4:0]    Axi4Incr_highCat;
  wire       [2:0]    Axi4Incr_sizeValue;
  wire       [11:0]   Axi4Incr_alignMask;
  wire       [11:0]   Axi4Incr_base;
  wire       [11:0]   Axi4Incr_baseIncr;
  reg        [1:0]    _zz_Axi4Incr_wrapCase;
  wire       [2:0]    Axi4Incr_wrapCase;
  wire                when_Axi4Channel_l307;
  wire                _zz_unburstify_result_ready;
  wire                stage0_valid;
  reg                 stage0_ready;
  wire                stage0_payload_last;
  wire       [16:0]   stage0_payload_fragment_addr;
  wire       [3:0]    stage0_payload_fragment_id;
  wire       [2:0]    stage0_payload_fragment_size;
  wire       [1:0]    stage0_payload_fragment_burst;
  wire                stage0_payload_fragment_write;
  wire       [14:0]   _zz_io_axi_r_payload_data;
  wire                stage0_fire;
  wire       [31:0]   _zz_io_axi_r_payload_data_1;
  wire                stage1_valid;
  wire                stage1_ready;
  wire                stage1_payload_last;
  wire       [16:0]   stage1_payload_fragment_addr;
  wire       [3:0]    stage1_payload_fragment_id;
  wire       [2:0]    stage1_payload_fragment_size;
  wire       [1:0]    stage1_payload_fragment_burst;
  wire                stage1_payload_fragment_write;
  reg                 stage0_rValid;
  reg                 stage0_rData_last;
  reg        [16:0]   stage0_rData_fragment_addr;
  reg        [3:0]    stage0_rData_fragment_id;
  reg        [2:0]    stage0_rData_fragment_size;
  reg        [1:0]    stage0_rData_fragment_burst;
  reg                 stage0_rData_fragment_write;
  wire                when_Stream_l368;
  reg [7:0] ram_symbol0 [0:32767];
  reg [7:0] ram_symbol1 [0:32767];
  reg [7:0] ram_symbol2 [0:32767];
  reg [7:0] ram_symbol3 [0:32767];
  reg [7:0] _zz_ramsymbol_read;
  reg [7:0] _zz_ramsymbol_read_1;
  reg [7:0] _zz_ramsymbol_read_2;
  reg [7:0] _zz_ramsymbol_read_3;

  assign _zz_Axi4Incr_alignMask = {(2'b01 < Axi4Incr_validSize),(2'b00 < Axi4Incr_validSize)};
  assign _zz_Axi4Incr_base_1 = unburstify_buffer_transaction_addr[11 : 0];
  assign _zz_Axi4Incr_base = _zz_Axi4Incr_base_1;
  assign _zz_Axi4Incr_baseIncr = {9'd0, Axi4Incr_sizeValue};
  assign _zz_Axi4Incr_wrapCase_1 = {1'd0, Axi4Incr_validSize};
  assign _zz_Axi4Incr_wrapCase_2 = {1'd0, _zz_Axi4Incr_wrapCase};
  assign _zz_Axi4Incr_result_1 = Axi4Incr_base[11 : 1];
  assign _zz_Axi4Incr_result_2 = Axi4Incr_baseIncr[0 : 0];
  assign _zz_Axi4Incr_result_3 = Axi4Incr_base[11 : 2];
  assign _zz_Axi4Incr_result_4 = Axi4Incr_baseIncr[1 : 0];
  assign _zz_Axi4Incr_result_5 = Axi4Incr_base[11 : 3];
  assign _zz_Axi4Incr_result_6 = Axi4Incr_baseIncr[2 : 0];
  assign _zz_Axi4Incr_result_7 = Axi4Incr_base[11 : 4];
  assign _zz_Axi4Incr_result_8 = Axi4Incr_baseIncr[3 : 0];
  assign _zz_Axi4Incr_result_9 = Axi4Incr_base[11 : 5];
  assign _zz_Axi4Incr_result_10 = Axi4Incr_baseIncr[4 : 0];
  assign _zz_Axi4Incr_result_11 = Axi4Incr_base[11 : 6];
  assign _zz_Axi4Incr_result_12 = Axi4Incr_baseIncr[5 : 0];
  initial begin
    $readmemb("DandSocSimple.v_toplevel_axi_bootram_ram_symbol0.bin",ram_symbol0);
    $readmemb("DandSocSimple.v_toplevel_axi_bootram_ram_symbol1.bin",ram_symbol1);
    $readmemb("DandSocSimple.v_toplevel_axi_bootram_ram_symbol2.bin",ram_symbol2);
    $readmemb("DandSocSimple.v_toplevel_axi_bootram_ram_symbol3.bin",ram_symbol3);
  end
  always @(*) begin
    _zz_ram_port0 = {_zz_ramsymbol_read_3, _zz_ramsymbol_read_2, _zz_ramsymbol_read_1, _zz_ramsymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(stage0_fire) begin
      _zz_ramsymbol_read <= ram_symbol0[_zz_io_axi_r_payload_data];
      _zz_ramsymbol_read_1 <= ram_symbol1[_zz_io_axi_r_payload_data];
      _zz_ramsymbol_read_2 <= ram_symbol2[_zz_io_axi_r_payload_data];
      _zz_ramsymbol_read_3 <= ram_symbol3[_zz_io_axi_r_payload_data];
    end
  end

  always @(posedge io_axiClk) begin
    if(io_axi_w_payload_strb[0] && stage0_fire && stage0_payload_fragment_write ) begin
      ram_symbol0[_zz_io_axi_r_payload_data] <= _zz_io_axi_r_payload_data_1[7 : 0];
    end
    if(io_axi_w_payload_strb[1] && stage0_fire && stage0_payload_fragment_write ) begin
      ram_symbol1[_zz_io_axi_r_payload_data] <= _zz_io_axi_r_payload_data_1[15 : 8];
    end
    if(io_axi_w_payload_strb[2] && stage0_fire && stage0_payload_fragment_write ) begin
      ram_symbol2[_zz_io_axi_r_payload_data] <= _zz_io_axi_r_payload_data_1[23 : 16];
    end
    if(io_axi_w_payload_strb[3] && stage0_fire && stage0_payload_fragment_write ) begin
      ram_symbol3[_zz_io_axi_r_payload_data] <= _zz_io_axi_r_payload_data_1[31 : 24];
    end
  end

  always @(*) begin
    case(Axi4Incr_wrapCase)
      3'b000 : _zz_Axi4Incr_result = {_zz_Axi4Incr_result_1,_zz_Axi4Incr_result_2};
      3'b001 : _zz_Axi4Incr_result = {_zz_Axi4Incr_result_3,_zz_Axi4Incr_result_4};
      3'b010 : _zz_Axi4Incr_result = {_zz_Axi4Incr_result_5,_zz_Axi4Incr_result_6};
      3'b011 : _zz_Axi4Incr_result = {_zz_Axi4Incr_result_7,_zz_Axi4Incr_result_8};
      3'b100 : _zz_Axi4Incr_result = {_zz_Axi4Incr_result_9,_zz_Axi4Incr_result_10};
      default : _zz_Axi4Incr_result = {_zz_Axi4Incr_result_11,_zz_Axi4Incr_result_12};
    endcase
  end

  assign unburstify_buffer_last = (unburstify_buffer_beat == 8'h01);
  assign Axi4Incr_validSize = unburstify_buffer_transaction_size[1 : 0];
  assign Axi4Incr_highCat = unburstify_buffer_transaction_addr[16 : 12];
  assign Axi4Incr_sizeValue = {(2'b10 == Axi4Incr_validSize),{(2'b01 == Axi4Incr_validSize),(2'b00 == Axi4Incr_validSize)}};
  assign Axi4Incr_alignMask = {10'd0, _zz_Axi4Incr_alignMask};
  assign Axi4Incr_base = (_zz_Axi4Incr_base & (~ Axi4Incr_alignMask));
  assign Axi4Incr_baseIncr = (Axi4Incr_base + _zz_Axi4Incr_baseIncr);
  always @(*) begin
    casez(unburstify_buffer_len)
      8'b????1??? : begin
        _zz_Axi4Incr_wrapCase = 2'b11;
      end
      8'b????01?? : begin
        _zz_Axi4Incr_wrapCase = 2'b10;
      end
      8'b????001? : begin
        _zz_Axi4Incr_wrapCase = 2'b01;
      end
      default : begin
        _zz_Axi4Incr_wrapCase = 2'b00;
      end
    endcase
  end

  assign Axi4Incr_wrapCase = (_zz_Axi4Incr_wrapCase_1 + _zz_Axi4Incr_wrapCase_2);
  always @(*) begin
    case(unburstify_buffer_transaction_burst)
      2'b00 : begin
        Axi4Incr_result = unburstify_buffer_transaction_addr;
      end
      2'b10 : begin
        Axi4Incr_result = {Axi4Incr_highCat,_zz_Axi4Incr_result};
      end
      default : begin
        Axi4Incr_result = {Axi4Incr_highCat,Axi4Incr_baseIncr};
      end
    endcase
  end

  always @(*) begin
    io_axi_arw_ready = 1'b0;
    if(!unburstify_buffer_valid) begin
      io_axi_arw_ready = unburstify_result_ready;
    end
  end

  always @(*) begin
    if(unburstify_buffer_valid) begin
      unburstify_result_valid = 1'b1;
    end else begin
      unburstify_result_valid = io_axi_arw_valid;
    end
  end

  always @(*) begin
    if(unburstify_buffer_valid) begin
      unburstify_result_payload_last = unburstify_buffer_last;
    end else begin
      unburstify_result_payload_last = 1'b1;
      if(when_Axi4Channel_l307) begin
        unburstify_result_payload_last = 1'b0;
      end
    end
  end

  always @(*) begin
    if(unburstify_buffer_valid) begin
      unburstify_result_payload_fragment_id = unburstify_buffer_transaction_id;
    end else begin
      unburstify_result_payload_fragment_id = io_axi_arw_payload_id;
    end
  end

  always @(*) begin
    if(unburstify_buffer_valid) begin
      unburstify_result_payload_fragment_size = unburstify_buffer_transaction_size;
    end else begin
      unburstify_result_payload_fragment_size = io_axi_arw_payload_size;
    end
  end

  always @(*) begin
    if(unburstify_buffer_valid) begin
      unburstify_result_payload_fragment_burst = unburstify_buffer_transaction_burst;
    end else begin
      unburstify_result_payload_fragment_burst = io_axi_arw_payload_burst;
    end
  end

  always @(*) begin
    if(unburstify_buffer_valid) begin
      unburstify_result_payload_fragment_write = unburstify_buffer_transaction_write;
    end else begin
      unburstify_result_payload_fragment_write = io_axi_arw_payload_write;
    end
  end

  always @(*) begin
    if(unburstify_buffer_valid) begin
      unburstify_result_payload_fragment_addr = Axi4Incr_result;
    end else begin
      unburstify_result_payload_fragment_addr = io_axi_arw_payload_addr;
    end
  end

  assign when_Axi4Channel_l307 = (io_axi_arw_payload_len != 8'h0);
  assign _zz_unburstify_result_ready = (! (unburstify_result_payload_fragment_write && (! io_axi_w_valid)));
  assign stage0_valid = (unburstify_result_valid && _zz_unburstify_result_ready);
  assign unburstify_result_ready = (stage0_ready && _zz_unburstify_result_ready);
  assign stage0_payload_last = unburstify_result_payload_last;
  assign stage0_payload_fragment_addr = unburstify_result_payload_fragment_addr;
  assign stage0_payload_fragment_id = unburstify_result_payload_fragment_id;
  assign stage0_payload_fragment_size = unburstify_result_payload_fragment_size;
  assign stage0_payload_fragment_burst = unburstify_result_payload_fragment_burst;
  assign stage0_payload_fragment_write = unburstify_result_payload_fragment_write;
  assign _zz_io_axi_r_payload_data = stage0_payload_fragment_addr[16 : 2];
  assign stage0_fire = (stage0_valid && stage0_ready);
  assign _zz_io_axi_r_payload_data_1 = io_axi_w_payload_data;
  assign io_axi_r_payload_data = _zz_ram_port0;
  assign io_axi_w_ready = ((unburstify_result_valid && unburstify_result_payload_fragment_write) && stage0_ready);
  always @(*) begin
    stage0_ready = stage1_ready;
    if(when_Stream_l368) begin
      stage0_ready = 1'b1;
    end
  end

  assign when_Stream_l368 = (! stage1_valid);
  assign stage1_valid = stage0_rValid;
  assign stage1_payload_last = stage0_rData_last;
  assign stage1_payload_fragment_addr = stage0_rData_fragment_addr;
  assign stage1_payload_fragment_id = stage0_rData_fragment_id;
  assign stage1_payload_fragment_size = stage0_rData_fragment_size;
  assign stage1_payload_fragment_burst = stage0_rData_fragment_burst;
  assign stage1_payload_fragment_write = stage0_rData_fragment_write;
  assign stage1_ready = ((io_axi_r_ready && (! stage1_payload_fragment_write)) || ((io_axi_b_ready || (! stage1_payload_last)) && stage1_payload_fragment_write));
  assign io_axi_r_valid = (stage1_valid && (! stage1_payload_fragment_write));
  assign io_axi_r_payload_id = stage1_payload_fragment_id;
  assign io_axi_r_payload_last = stage1_payload_last;
  assign io_axi_r_payload_resp = 2'b00;
  assign io_axi_b_valid = ((stage1_valid && stage1_payload_fragment_write) && stage1_payload_last);
  assign io_axi_b_payload_resp = 2'b00;
  assign io_axi_b_payload_id = stage1_payload_fragment_id;
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      unburstify_buffer_valid <= 1'b0;
      stage0_rValid <= 1'b0;
    end else begin
      if(unburstify_result_ready) begin
        if(unburstify_buffer_last) begin
          unburstify_buffer_valid <= 1'b0;
        end
      end
      if(!unburstify_buffer_valid) begin
        if(when_Axi4Channel_l307) begin
          if(unburstify_result_ready) begin
            unburstify_buffer_valid <= io_axi_arw_valid;
          end
        end
      end
      if(stage0_ready) begin
        stage0_rValid <= stage0_valid;
      end
    end
  end

  always @(posedge io_axiClk) begin
    if(unburstify_result_ready) begin
      unburstify_buffer_beat <= (unburstify_buffer_beat - 8'h01);
      unburstify_buffer_transaction_addr[11 : 0] <= Axi4Incr_result[11 : 0];
    end
    if(!unburstify_buffer_valid) begin
      if(when_Axi4Channel_l307) begin
        if(unburstify_result_ready) begin
          unburstify_buffer_transaction_addr <= io_axi_arw_payload_addr;
          unburstify_buffer_transaction_id <= io_axi_arw_payload_id;
          unburstify_buffer_transaction_size <= io_axi_arw_payload_size;
          unburstify_buffer_transaction_burst <= io_axi_arw_payload_burst;
          unburstify_buffer_transaction_write <= io_axi_arw_payload_write;
          unburstify_buffer_beat <= io_axi_arw_payload_len;
          unburstify_buffer_len <= io_axi_arw_payload_len;
        end
      end
    end
    if(stage0_ready) begin
      stage0_rData_last <= stage0_payload_last;
      stage0_rData_fragment_addr <= stage0_payload_fragment_addr;
      stage0_rData_fragment_id <= stage0_payload_fragment_id;
      stage0_rData_fragment_size <= stage0_payload_fragment_size;
      stage0_rData_fragment_burst <= stage0_payload_fragment_burst;
      stage0_rData_fragment_write <= stage0_payload_fragment_write;
    end
  end


endmodule

module Axi4SharedOnChipRam (
  input               io_axi_arw_valid,
  output reg          io_axi_arw_ready,
  input      [16:0]   io_axi_arw_payload_addr,
  input      [3:0]    io_axi_arw_payload_id,
  input      [7:0]    io_axi_arw_payload_len,
  input      [2:0]    io_axi_arw_payload_size,
  input      [1:0]    io_axi_arw_payload_burst,
  input               io_axi_arw_payload_write,
  input               io_axi_w_valid,
  output              io_axi_w_ready,
  input      [63:0]   io_axi_w_payload_data,
  input      [7:0]    io_axi_w_payload_strb,
  input               io_axi_w_payload_last,
  output              io_axi_b_valid,
  input               io_axi_b_ready,
  output     [3:0]    io_axi_b_payload_id,
  output     [1:0]    io_axi_b_payload_resp,
  output              io_axi_r_valid,
  input               io_axi_r_ready,
  output     [63:0]   io_axi_r_payload_data,
  output     [3:0]    io_axi_r_payload_id,
  output     [1:0]    io_axi_r_payload_resp,
  output              io_axi_r_payload_last,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  reg        [63:0]   _zz_ram_port0;
  wire       [2:0]    _zz_Axi4Incr_alignMask;
  wire       [11:0]   _zz_Axi4Incr_base;
  wire       [11:0]   _zz_Axi4Incr_base_1;
  wire       [11:0]   _zz_Axi4Incr_baseIncr;
  wire       [2:0]    _zz_Axi4Incr_wrapCase_1;
  wire       [2:0]    _zz_Axi4Incr_wrapCase_2;
  reg        [11:0]   _zz_Axi4Incr_result;
  wire       [10:0]   _zz_Axi4Incr_result_1;
  wire       [0:0]    _zz_Axi4Incr_result_2;
  wire       [9:0]    _zz_Axi4Incr_result_3;
  wire       [1:0]    _zz_Axi4Incr_result_4;
  wire       [8:0]    _zz_Axi4Incr_result_5;
  wire       [2:0]    _zz_Axi4Incr_result_6;
  wire       [7:0]    _zz_Axi4Incr_result_7;
  wire       [3:0]    _zz_Axi4Incr_result_8;
  wire       [6:0]    _zz_Axi4Incr_result_9;
  wire       [4:0]    _zz_Axi4Incr_result_10;
  wire       [5:0]    _zz_Axi4Incr_result_11;
  wire       [5:0]    _zz_Axi4Incr_result_12;
  wire       [4:0]    _zz_Axi4Incr_result_13;
  wire       [6:0]    _zz_Axi4Incr_result_14;
  reg                 unburstify_result_valid;
  wire                unburstify_result_ready;
  reg                 unburstify_result_payload_last;
  reg        [16:0]   unburstify_result_payload_fragment_addr;
  reg        [3:0]    unburstify_result_payload_fragment_id;
  reg        [2:0]    unburstify_result_payload_fragment_size;
  reg        [1:0]    unburstify_result_payload_fragment_burst;
  reg                 unburstify_result_payload_fragment_write;
  wire                unburstify_doResult;
  reg                 unburstify_buffer_valid;
  reg        [7:0]    unburstify_buffer_len;
  reg        [7:0]    unburstify_buffer_beat;
  reg        [16:0]   unburstify_buffer_transaction_addr;
  reg        [3:0]    unburstify_buffer_transaction_id;
  reg        [2:0]    unburstify_buffer_transaction_size;
  reg        [1:0]    unburstify_buffer_transaction_burst;
  reg                 unburstify_buffer_transaction_write;
  wire                unburstify_buffer_last;
  wire       [1:0]    Axi4Incr_validSize;
  reg        [16:0]   Axi4Incr_result;
  wire       [4:0]    Axi4Incr_highCat;
  wire       [3:0]    Axi4Incr_sizeValue;
  wire       [11:0]   Axi4Incr_alignMask;
  wire       [11:0]   Axi4Incr_base;
  wire       [11:0]   Axi4Incr_baseIncr;
  reg        [1:0]    _zz_Axi4Incr_wrapCase;
  wire       [2:0]    Axi4Incr_wrapCase;
  wire                when_Axi4Channel_l307;
  wire                _zz_unburstify_result_ready;
  wire                stage0_valid;
  reg                 stage0_ready;
  wire                stage0_payload_last;
  wire       [16:0]   stage0_payload_fragment_addr;
  wire       [3:0]    stage0_payload_fragment_id;
  wire       [2:0]    stage0_payload_fragment_size;
  wire       [1:0]    stage0_payload_fragment_burst;
  wire                stage0_payload_fragment_write;
  wire       [13:0]   _zz_io_axi_r_payload_data;
  wire                stage0_fire;
  wire       [63:0]   _zz_io_axi_r_payload_data_1;
  wire                stage1_valid;
  wire                stage1_ready;
  wire                stage1_payload_last;
  wire       [16:0]   stage1_payload_fragment_addr;
  wire       [3:0]    stage1_payload_fragment_id;
  wire       [2:0]    stage1_payload_fragment_size;
  wire       [1:0]    stage1_payload_fragment_burst;
  wire                stage1_payload_fragment_write;
  reg                 stage0_rValid;
  reg                 stage0_rData_last;
  reg        [16:0]   stage0_rData_fragment_addr;
  reg        [3:0]    stage0_rData_fragment_id;
  reg        [2:0]    stage0_rData_fragment_size;
  reg        [1:0]    stage0_rData_fragment_burst;
  reg                 stage0_rData_fragment_write;
  wire                when_Stream_l368;
  reg [7:0] ram_symbol0 [0:16383];
  reg [7:0] ram_symbol1 [0:16383];
  reg [7:0] ram_symbol2 [0:16383];
  reg [7:0] ram_symbol3 [0:16383];
  reg [7:0] ram_symbol4 [0:16383];
  reg [7:0] ram_symbol5 [0:16383];
  reg [7:0] ram_symbol6 [0:16383];
  reg [7:0] ram_symbol7 [0:16383];
  reg [7:0] _zz_ramsymbol_read;
  reg [7:0] _zz_ramsymbol_read_1;
  reg [7:0] _zz_ramsymbol_read_2;
  reg [7:0] _zz_ramsymbol_read_3;
  reg [7:0] _zz_ramsymbol_read_4;
  reg [7:0] _zz_ramsymbol_read_5;
  reg [7:0] _zz_ramsymbol_read_6;
  reg [7:0] _zz_ramsymbol_read_7;

  assign _zz_Axi4Incr_alignMask = {(2'b10 < Axi4Incr_validSize),{(2'b01 < Axi4Incr_validSize),(2'b00 < Axi4Incr_validSize)}};
  assign _zz_Axi4Incr_base_1 = unburstify_buffer_transaction_addr[11 : 0];
  assign _zz_Axi4Incr_base = _zz_Axi4Incr_base_1;
  assign _zz_Axi4Incr_baseIncr = {8'd0, Axi4Incr_sizeValue};
  assign _zz_Axi4Incr_wrapCase_1 = {1'd0, Axi4Incr_validSize};
  assign _zz_Axi4Incr_wrapCase_2 = {1'd0, _zz_Axi4Incr_wrapCase};
  assign _zz_Axi4Incr_result_1 = Axi4Incr_base[11 : 1];
  assign _zz_Axi4Incr_result_2 = Axi4Incr_baseIncr[0 : 0];
  assign _zz_Axi4Incr_result_3 = Axi4Incr_base[11 : 2];
  assign _zz_Axi4Incr_result_4 = Axi4Incr_baseIncr[1 : 0];
  assign _zz_Axi4Incr_result_5 = Axi4Incr_base[11 : 3];
  assign _zz_Axi4Incr_result_6 = Axi4Incr_baseIncr[2 : 0];
  assign _zz_Axi4Incr_result_7 = Axi4Incr_base[11 : 4];
  assign _zz_Axi4Incr_result_8 = Axi4Incr_baseIncr[3 : 0];
  assign _zz_Axi4Incr_result_9 = Axi4Incr_base[11 : 5];
  assign _zz_Axi4Incr_result_10 = Axi4Incr_baseIncr[4 : 0];
  assign _zz_Axi4Incr_result_11 = Axi4Incr_base[11 : 6];
  assign _zz_Axi4Incr_result_12 = Axi4Incr_baseIncr[5 : 0];
  assign _zz_Axi4Incr_result_13 = Axi4Incr_base[11 : 7];
  assign _zz_Axi4Incr_result_14 = Axi4Incr_baseIncr[6 : 0];
  always @(*) begin
    _zz_ram_port0 = {_zz_ramsymbol_read_7, _zz_ramsymbol_read_6, _zz_ramsymbol_read_5, _zz_ramsymbol_read_4, _zz_ramsymbol_read_3, _zz_ramsymbol_read_2, _zz_ramsymbol_read_1, _zz_ramsymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(stage0_fire) begin
      _zz_ramsymbol_read <= ram_symbol0[_zz_io_axi_r_payload_data];
      _zz_ramsymbol_read_1 <= ram_symbol1[_zz_io_axi_r_payload_data];
      _zz_ramsymbol_read_2 <= ram_symbol2[_zz_io_axi_r_payload_data];
      _zz_ramsymbol_read_3 <= ram_symbol3[_zz_io_axi_r_payload_data];
      _zz_ramsymbol_read_4 <= ram_symbol4[_zz_io_axi_r_payload_data];
      _zz_ramsymbol_read_5 <= ram_symbol5[_zz_io_axi_r_payload_data];
      _zz_ramsymbol_read_6 <= ram_symbol6[_zz_io_axi_r_payload_data];
      _zz_ramsymbol_read_7 <= ram_symbol7[_zz_io_axi_r_payload_data];
    end
  end

  always @(posedge io_axiClk) begin
    if(io_axi_w_payload_strb[0] && stage0_fire && stage0_payload_fragment_write ) begin
      ram_symbol0[_zz_io_axi_r_payload_data] <= _zz_io_axi_r_payload_data_1[7 : 0];
    end
    if(io_axi_w_payload_strb[1] && stage0_fire && stage0_payload_fragment_write ) begin
      ram_symbol1[_zz_io_axi_r_payload_data] <= _zz_io_axi_r_payload_data_1[15 : 8];
    end
    if(io_axi_w_payload_strb[2] && stage0_fire && stage0_payload_fragment_write ) begin
      ram_symbol2[_zz_io_axi_r_payload_data] <= _zz_io_axi_r_payload_data_1[23 : 16];
    end
    if(io_axi_w_payload_strb[3] && stage0_fire && stage0_payload_fragment_write ) begin
      ram_symbol3[_zz_io_axi_r_payload_data] <= _zz_io_axi_r_payload_data_1[31 : 24];
    end
    if(io_axi_w_payload_strb[4] && stage0_fire && stage0_payload_fragment_write ) begin
      ram_symbol4[_zz_io_axi_r_payload_data] <= _zz_io_axi_r_payload_data_1[39 : 32];
    end
    if(io_axi_w_payload_strb[5] && stage0_fire && stage0_payload_fragment_write ) begin
      ram_symbol5[_zz_io_axi_r_payload_data] <= _zz_io_axi_r_payload_data_1[47 : 40];
    end
    if(io_axi_w_payload_strb[6] && stage0_fire && stage0_payload_fragment_write ) begin
      ram_symbol6[_zz_io_axi_r_payload_data] <= _zz_io_axi_r_payload_data_1[55 : 48];
    end
    if(io_axi_w_payload_strb[7] && stage0_fire && stage0_payload_fragment_write ) begin
      ram_symbol7[_zz_io_axi_r_payload_data] <= _zz_io_axi_r_payload_data_1[63 : 56];
    end
  end

  always @(*) begin
    case(Axi4Incr_wrapCase)
      3'b000 : _zz_Axi4Incr_result = {_zz_Axi4Incr_result_1,_zz_Axi4Incr_result_2};
      3'b001 : _zz_Axi4Incr_result = {_zz_Axi4Incr_result_3,_zz_Axi4Incr_result_4};
      3'b010 : _zz_Axi4Incr_result = {_zz_Axi4Incr_result_5,_zz_Axi4Incr_result_6};
      3'b011 : _zz_Axi4Incr_result = {_zz_Axi4Incr_result_7,_zz_Axi4Incr_result_8};
      3'b100 : _zz_Axi4Incr_result = {_zz_Axi4Incr_result_9,_zz_Axi4Incr_result_10};
      3'b101 : _zz_Axi4Incr_result = {_zz_Axi4Incr_result_11,_zz_Axi4Incr_result_12};
      default : _zz_Axi4Incr_result = {_zz_Axi4Incr_result_13,_zz_Axi4Incr_result_14};
    endcase
  end

  assign unburstify_buffer_last = (unburstify_buffer_beat == 8'h01);
  assign Axi4Incr_validSize = unburstify_buffer_transaction_size[1 : 0];
  assign Axi4Incr_highCat = unburstify_buffer_transaction_addr[16 : 12];
  assign Axi4Incr_sizeValue = {(2'b11 == Axi4Incr_validSize),{(2'b10 == Axi4Incr_validSize),{(2'b01 == Axi4Incr_validSize),(2'b00 == Axi4Incr_validSize)}}};
  assign Axi4Incr_alignMask = {9'd0, _zz_Axi4Incr_alignMask};
  assign Axi4Incr_base = (_zz_Axi4Incr_base & (~ Axi4Incr_alignMask));
  assign Axi4Incr_baseIncr = (Axi4Incr_base + _zz_Axi4Incr_baseIncr);
  always @(*) begin
    casez(unburstify_buffer_len)
      8'b????1??? : begin
        _zz_Axi4Incr_wrapCase = 2'b11;
      end
      8'b????01?? : begin
        _zz_Axi4Incr_wrapCase = 2'b10;
      end
      8'b????001? : begin
        _zz_Axi4Incr_wrapCase = 2'b01;
      end
      default : begin
        _zz_Axi4Incr_wrapCase = 2'b00;
      end
    endcase
  end

  assign Axi4Incr_wrapCase = (_zz_Axi4Incr_wrapCase_1 + _zz_Axi4Incr_wrapCase_2);
  always @(*) begin
    case(unburstify_buffer_transaction_burst)
      2'b00 : begin
        Axi4Incr_result = unburstify_buffer_transaction_addr;
      end
      2'b10 : begin
        Axi4Incr_result = {Axi4Incr_highCat,_zz_Axi4Incr_result};
      end
      default : begin
        Axi4Incr_result = {Axi4Incr_highCat,Axi4Incr_baseIncr};
      end
    endcase
  end

  always @(*) begin
    io_axi_arw_ready = 1'b0;
    if(!unburstify_buffer_valid) begin
      io_axi_arw_ready = unburstify_result_ready;
    end
  end

  always @(*) begin
    if(unburstify_buffer_valid) begin
      unburstify_result_valid = 1'b1;
    end else begin
      unburstify_result_valid = io_axi_arw_valid;
    end
  end

  always @(*) begin
    if(unburstify_buffer_valid) begin
      unburstify_result_payload_last = unburstify_buffer_last;
    end else begin
      unburstify_result_payload_last = 1'b1;
      if(when_Axi4Channel_l307) begin
        unburstify_result_payload_last = 1'b0;
      end
    end
  end

  always @(*) begin
    if(unburstify_buffer_valid) begin
      unburstify_result_payload_fragment_id = unburstify_buffer_transaction_id;
    end else begin
      unburstify_result_payload_fragment_id = io_axi_arw_payload_id;
    end
  end

  always @(*) begin
    if(unburstify_buffer_valid) begin
      unburstify_result_payload_fragment_size = unburstify_buffer_transaction_size;
    end else begin
      unburstify_result_payload_fragment_size = io_axi_arw_payload_size;
    end
  end

  always @(*) begin
    if(unburstify_buffer_valid) begin
      unburstify_result_payload_fragment_burst = unburstify_buffer_transaction_burst;
    end else begin
      unburstify_result_payload_fragment_burst = io_axi_arw_payload_burst;
    end
  end

  always @(*) begin
    if(unburstify_buffer_valid) begin
      unburstify_result_payload_fragment_write = unburstify_buffer_transaction_write;
    end else begin
      unburstify_result_payload_fragment_write = io_axi_arw_payload_write;
    end
  end

  always @(*) begin
    if(unburstify_buffer_valid) begin
      unburstify_result_payload_fragment_addr = Axi4Incr_result;
    end else begin
      unburstify_result_payload_fragment_addr = io_axi_arw_payload_addr;
    end
  end

  assign when_Axi4Channel_l307 = (io_axi_arw_payload_len != 8'h0);
  assign _zz_unburstify_result_ready = (! (unburstify_result_payload_fragment_write && (! io_axi_w_valid)));
  assign stage0_valid = (unburstify_result_valid && _zz_unburstify_result_ready);
  assign unburstify_result_ready = (stage0_ready && _zz_unburstify_result_ready);
  assign stage0_payload_last = unburstify_result_payload_last;
  assign stage0_payload_fragment_addr = unburstify_result_payload_fragment_addr;
  assign stage0_payload_fragment_id = unburstify_result_payload_fragment_id;
  assign stage0_payload_fragment_size = unburstify_result_payload_fragment_size;
  assign stage0_payload_fragment_burst = unburstify_result_payload_fragment_burst;
  assign stage0_payload_fragment_write = unburstify_result_payload_fragment_write;
  assign _zz_io_axi_r_payload_data = stage0_payload_fragment_addr[16 : 3];
  assign stage0_fire = (stage0_valid && stage0_ready);
  assign _zz_io_axi_r_payload_data_1 = io_axi_w_payload_data;
  assign io_axi_r_payload_data = _zz_ram_port0;
  assign io_axi_w_ready = ((unburstify_result_valid && unburstify_result_payload_fragment_write) && stage0_ready);
  always @(*) begin
    stage0_ready = stage1_ready;
    if(when_Stream_l368) begin
      stage0_ready = 1'b1;
    end
  end

  assign when_Stream_l368 = (! stage1_valid);
  assign stage1_valid = stage0_rValid;
  assign stage1_payload_last = stage0_rData_last;
  assign stage1_payload_fragment_addr = stage0_rData_fragment_addr;
  assign stage1_payload_fragment_id = stage0_rData_fragment_id;
  assign stage1_payload_fragment_size = stage0_rData_fragment_size;
  assign stage1_payload_fragment_burst = stage0_rData_fragment_burst;
  assign stage1_payload_fragment_write = stage0_rData_fragment_write;
  assign stage1_ready = ((io_axi_r_ready && (! stage1_payload_fragment_write)) || ((io_axi_b_ready || (! stage1_payload_last)) && stage1_payload_fragment_write));
  assign io_axi_r_valid = (stage1_valid && (! stage1_payload_fragment_write));
  assign io_axi_r_payload_id = stage1_payload_fragment_id;
  assign io_axi_r_payload_last = stage1_payload_last;
  assign io_axi_r_payload_resp = 2'b00;
  assign io_axi_b_valid = ((stage1_valid && stage1_payload_fragment_write) && stage1_payload_last);
  assign io_axi_b_payload_resp = 2'b00;
  assign io_axi_b_payload_id = stage1_payload_fragment_id;
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      unburstify_buffer_valid <= 1'b0;
      stage0_rValid <= 1'b0;
    end else begin
      if(unburstify_result_ready) begin
        if(unburstify_buffer_last) begin
          unburstify_buffer_valid <= 1'b0;
        end
      end
      if(!unburstify_buffer_valid) begin
        if(when_Axi4Channel_l307) begin
          if(unburstify_result_ready) begin
            unburstify_buffer_valid <= io_axi_arw_valid;
          end
        end
      end
      if(stage0_ready) begin
        stage0_rValid <= stage0_valid;
      end
    end
  end

  always @(posedge io_axiClk) begin
    if(unburstify_result_ready) begin
      unburstify_buffer_beat <= (unburstify_buffer_beat - 8'h01);
      unburstify_buffer_transaction_addr[11 : 0] <= Axi4Incr_result[11 : 0];
    end
    if(!unburstify_buffer_valid) begin
      if(when_Axi4Channel_l307) begin
        if(unburstify_result_ready) begin
          unburstify_buffer_transaction_addr <= io_axi_arw_payload_addr;
          unburstify_buffer_transaction_id <= io_axi_arw_payload_id;
          unburstify_buffer_transaction_size <= io_axi_arw_payload_size;
          unburstify_buffer_transaction_burst <= io_axi_arw_payload_burst;
          unburstify_buffer_transaction_write <= io_axi_arw_payload_write;
          unburstify_buffer_beat <= io_axi_arw_payload_len;
          unburstify_buffer_len <= io_axi_arw_payload_len;
        end
      end
    end
    if(stage0_ready) begin
      stage0_rData_last <= stage0_payload_last;
      stage0_rData_fragment_addr <= stage0_payload_fragment_addr;
      stage0_rData_fragment_id <= stage0_payload_fragment_id;
      stage0_rData_fragment_size <= stage0_payload_fragment_size;
      stage0_rData_fragment_burst <= stage0_payload_fragment_burst;
      stage0_rData_fragment_write <= stage0_payload_fragment_write;
    end
  end


endmodule

module Axi4Downsizer (
  input               io_input_aw_valid,
  output              io_input_aw_ready,
  input      [31:0]   io_input_aw_payload_addr,
  input      [3:0]    io_input_aw_payload_id,
  input      [3:0]    io_input_aw_payload_region,
  input      [7:0]    io_input_aw_payload_len,
  input      [2:0]    io_input_aw_payload_size,
  input      [1:0]    io_input_aw_payload_burst,
  input      [0:0]    io_input_aw_payload_lock,
  input      [3:0]    io_input_aw_payload_cache,
  input      [3:0]    io_input_aw_payload_qos,
  input      [2:0]    io_input_aw_payload_prot,
  input               io_input_w_valid,
  output              io_input_w_ready,
  input      [63:0]   io_input_w_payload_data,
  input      [7:0]    io_input_w_payload_strb,
  input               io_input_w_payload_last,
  output              io_input_b_valid,
  input               io_input_b_ready,
  output     [3:0]    io_input_b_payload_id,
  output     [1:0]    io_input_b_payload_resp,
  input               io_input_ar_valid,
  output              io_input_ar_ready,
  input      [31:0]   io_input_ar_payload_addr,
  input      [3:0]    io_input_ar_payload_id,
  input      [3:0]    io_input_ar_payload_region,
  input      [7:0]    io_input_ar_payload_len,
  input      [2:0]    io_input_ar_payload_size,
  input      [1:0]    io_input_ar_payload_burst,
  input      [0:0]    io_input_ar_payload_lock,
  input      [3:0]    io_input_ar_payload_cache,
  input      [3:0]    io_input_ar_payload_qos,
  input      [2:0]    io_input_ar_payload_prot,
  output              io_input_r_valid,
  input               io_input_r_ready,
  output     [63:0]   io_input_r_payload_data,
  output     [3:0]    io_input_r_payload_id,
  output     [1:0]    io_input_r_payload_resp,
  output              io_input_r_payload_last,
  output              io_output_aw_valid,
  input               io_output_aw_ready,
  output     [31:0]   io_output_aw_payload_addr,
  output     [3:0]    io_output_aw_payload_id,
  output     [3:0]    io_output_aw_payload_region,
  output     [7:0]    io_output_aw_payload_len,
  output     [2:0]    io_output_aw_payload_size,
  output     [1:0]    io_output_aw_payload_burst,
  output     [0:0]    io_output_aw_payload_lock,
  output     [3:0]    io_output_aw_payload_cache,
  output     [3:0]    io_output_aw_payload_qos,
  output     [2:0]    io_output_aw_payload_prot,
  output              io_output_w_valid,
  input               io_output_w_ready,
  output     [31:0]   io_output_w_payload_data,
  output     [3:0]    io_output_w_payload_strb,
  output              io_output_w_payload_last,
  input               io_output_b_valid,
  output              io_output_b_ready,
  input      [3:0]    io_output_b_payload_id,
  input      [1:0]    io_output_b_payload_resp,
  output              io_output_ar_valid,
  input               io_output_ar_ready,
  output     [31:0]   io_output_ar_payload_addr,
  output     [3:0]    io_output_ar_payload_id,
  output     [3:0]    io_output_ar_payload_region,
  output     [7:0]    io_output_ar_payload_len,
  output     [2:0]    io_output_ar_payload_size,
  output     [1:0]    io_output_ar_payload_burst,
  output     [0:0]    io_output_ar_payload_lock,
  output     [3:0]    io_output_ar_payload_cache,
  output     [3:0]    io_output_ar_payload_qos,
  output     [2:0]    io_output_ar_payload_prot,
  input               io_output_r_valid,
  output              io_output_r_ready,
  input      [31:0]   io_output_r_payload_data,
  input      [3:0]    io_output_r_payload_id,
  input      [1:0]    io_output_r_payload_resp,
  input               io_output_r_payload_last,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  wire                readOnly_io_input_ar_ready;
  wire                readOnly_io_input_r_valid;
  wire       [63:0]   readOnly_io_input_r_payload_data;
  wire       [3:0]    readOnly_io_input_r_payload_id;
  wire       [1:0]    readOnly_io_input_r_payload_resp;
  wire                readOnly_io_input_r_payload_last;
  wire                readOnly_io_output_ar_valid;
  wire       [31:0]   readOnly_io_output_ar_payload_addr;
  wire       [3:0]    readOnly_io_output_ar_payload_id;
  wire       [3:0]    readOnly_io_output_ar_payload_region;
  wire       [7:0]    readOnly_io_output_ar_payload_len;
  wire       [2:0]    readOnly_io_output_ar_payload_size;
  wire       [1:0]    readOnly_io_output_ar_payload_burst;
  wire       [0:0]    readOnly_io_output_ar_payload_lock;
  wire       [3:0]    readOnly_io_output_ar_payload_cache;
  wire       [3:0]    readOnly_io_output_ar_payload_qos;
  wire       [2:0]    readOnly_io_output_ar_payload_prot;
  wire                readOnly_io_output_r_ready;
  wire                writeOnly_io_input_aw_ready;
  wire                writeOnly_io_input_w_ready;
  wire                writeOnly_io_input_b_valid;
  wire       [3:0]    writeOnly_io_input_b_payload_id;
  wire       [1:0]    writeOnly_io_input_b_payload_resp;
  wire                writeOnly_io_output_aw_valid;
  wire       [31:0]   writeOnly_io_output_aw_payload_addr;
  wire       [3:0]    writeOnly_io_output_aw_payload_id;
  wire       [3:0]    writeOnly_io_output_aw_payload_region;
  wire       [7:0]    writeOnly_io_output_aw_payload_len;
  wire       [2:0]    writeOnly_io_output_aw_payload_size;
  wire       [1:0]    writeOnly_io_output_aw_payload_burst;
  wire       [0:0]    writeOnly_io_output_aw_payload_lock;
  wire       [3:0]    writeOnly_io_output_aw_payload_cache;
  wire       [3:0]    writeOnly_io_output_aw_payload_qos;
  wire       [2:0]    writeOnly_io_output_aw_payload_prot;
  wire                writeOnly_io_output_w_valid;
  wire       [31:0]   writeOnly_io_output_w_payload_data;
  wire       [3:0]    writeOnly_io_output_w_payload_strb;
  wire                writeOnly_io_output_w_payload_last;
  wire                writeOnly_io_output_b_ready;

  Axi4ReadOnlyDownsizer readOnly (
    .io_input_ar_valid           (io_input_ar_valid                        ), //i
    .io_input_ar_ready           (readOnly_io_input_ar_ready               ), //o
    .io_input_ar_payload_addr    (io_input_ar_payload_addr[31:0]           ), //i
    .io_input_ar_payload_id      (io_input_ar_payload_id[3:0]              ), //i
    .io_input_ar_payload_region  (io_input_ar_payload_region[3:0]          ), //i
    .io_input_ar_payload_len     (io_input_ar_payload_len[7:0]             ), //i
    .io_input_ar_payload_size    (io_input_ar_payload_size[2:0]            ), //i
    .io_input_ar_payload_burst   (io_input_ar_payload_burst[1:0]           ), //i
    .io_input_ar_payload_lock    (io_input_ar_payload_lock                 ), //i
    .io_input_ar_payload_cache   (io_input_ar_payload_cache[3:0]           ), //i
    .io_input_ar_payload_qos     (io_input_ar_payload_qos[3:0]             ), //i
    .io_input_ar_payload_prot    (io_input_ar_payload_prot[2:0]            ), //i
    .io_input_r_valid            (readOnly_io_input_r_valid                ), //o
    .io_input_r_ready            (io_input_r_ready                         ), //i
    .io_input_r_payload_data     (readOnly_io_input_r_payload_data[63:0]   ), //o
    .io_input_r_payload_id       (readOnly_io_input_r_payload_id[3:0]      ), //o
    .io_input_r_payload_resp     (readOnly_io_input_r_payload_resp[1:0]    ), //o
    .io_input_r_payload_last     (readOnly_io_input_r_payload_last         ), //o
    .io_output_ar_valid          (readOnly_io_output_ar_valid              ), //o
    .io_output_ar_ready          (io_output_ar_ready                       ), //i
    .io_output_ar_payload_addr   (readOnly_io_output_ar_payload_addr[31:0] ), //o
    .io_output_ar_payload_id     (readOnly_io_output_ar_payload_id[3:0]    ), //o
    .io_output_ar_payload_region (readOnly_io_output_ar_payload_region[3:0]), //o
    .io_output_ar_payload_len    (readOnly_io_output_ar_payload_len[7:0]   ), //o
    .io_output_ar_payload_size   (readOnly_io_output_ar_payload_size[2:0]  ), //o
    .io_output_ar_payload_burst  (readOnly_io_output_ar_payload_burst[1:0] ), //o
    .io_output_ar_payload_lock   (readOnly_io_output_ar_payload_lock       ), //o
    .io_output_ar_payload_cache  (readOnly_io_output_ar_payload_cache[3:0] ), //o
    .io_output_ar_payload_qos    (readOnly_io_output_ar_payload_qos[3:0]   ), //o
    .io_output_ar_payload_prot   (readOnly_io_output_ar_payload_prot[2:0]  ), //o
    .io_output_r_valid           (io_output_r_valid                        ), //i
    .io_output_r_ready           (readOnly_io_output_r_ready               ), //o
    .io_output_r_payload_data    (io_output_r_payload_data[31:0]           ), //i
    .io_output_r_payload_id      (io_output_r_payload_id[3:0]              ), //i
    .io_output_r_payload_resp    (io_output_r_payload_resp[1:0]            ), //i
    .io_output_r_payload_last    (io_output_r_payload_last                 ), //i
    .io_axiClk                   (io_axiClk                                ), //i
    .resetCtrl_axiReset          (resetCtrl_axiReset                       )  //i
  );
  Axi4WriteOnlyDownsizer writeOnly (
    .io_input_aw_valid           (io_input_aw_valid                         ), //i
    .io_input_aw_ready           (writeOnly_io_input_aw_ready               ), //o
    .io_input_aw_payload_addr    (io_input_aw_payload_addr[31:0]            ), //i
    .io_input_aw_payload_id      (io_input_aw_payload_id[3:0]               ), //i
    .io_input_aw_payload_region  (io_input_aw_payload_region[3:0]           ), //i
    .io_input_aw_payload_len     (io_input_aw_payload_len[7:0]              ), //i
    .io_input_aw_payload_size    (io_input_aw_payload_size[2:0]             ), //i
    .io_input_aw_payload_burst   (io_input_aw_payload_burst[1:0]            ), //i
    .io_input_aw_payload_lock    (io_input_aw_payload_lock                  ), //i
    .io_input_aw_payload_cache   (io_input_aw_payload_cache[3:0]            ), //i
    .io_input_aw_payload_qos     (io_input_aw_payload_qos[3:0]              ), //i
    .io_input_aw_payload_prot    (io_input_aw_payload_prot[2:0]             ), //i
    .io_input_w_valid            (io_input_w_valid                          ), //i
    .io_input_w_ready            (writeOnly_io_input_w_ready                ), //o
    .io_input_w_payload_data     (io_input_w_payload_data[63:0]             ), //i
    .io_input_w_payload_strb     (io_input_w_payload_strb[7:0]              ), //i
    .io_input_w_payload_last     (io_input_w_payload_last                   ), //i
    .io_input_b_valid            (writeOnly_io_input_b_valid                ), //o
    .io_input_b_ready            (io_input_b_ready                          ), //i
    .io_input_b_payload_id       (writeOnly_io_input_b_payload_id[3:0]      ), //o
    .io_input_b_payload_resp     (writeOnly_io_input_b_payload_resp[1:0]    ), //o
    .io_output_aw_valid          (writeOnly_io_output_aw_valid              ), //o
    .io_output_aw_ready          (io_output_aw_ready                        ), //i
    .io_output_aw_payload_addr   (writeOnly_io_output_aw_payload_addr[31:0] ), //o
    .io_output_aw_payload_id     (writeOnly_io_output_aw_payload_id[3:0]    ), //o
    .io_output_aw_payload_region (writeOnly_io_output_aw_payload_region[3:0]), //o
    .io_output_aw_payload_len    (writeOnly_io_output_aw_payload_len[7:0]   ), //o
    .io_output_aw_payload_size   (writeOnly_io_output_aw_payload_size[2:0]  ), //o
    .io_output_aw_payload_burst  (writeOnly_io_output_aw_payload_burst[1:0] ), //o
    .io_output_aw_payload_lock   (writeOnly_io_output_aw_payload_lock       ), //o
    .io_output_aw_payload_cache  (writeOnly_io_output_aw_payload_cache[3:0] ), //o
    .io_output_aw_payload_qos    (writeOnly_io_output_aw_payload_qos[3:0]   ), //o
    .io_output_aw_payload_prot   (writeOnly_io_output_aw_payload_prot[2:0]  ), //o
    .io_output_w_valid           (writeOnly_io_output_w_valid               ), //o
    .io_output_w_ready           (io_output_w_ready                         ), //i
    .io_output_w_payload_data    (writeOnly_io_output_w_payload_data[31:0]  ), //o
    .io_output_w_payload_strb    (writeOnly_io_output_w_payload_strb[3:0]   ), //o
    .io_output_w_payload_last    (writeOnly_io_output_w_payload_last        ), //o
    .io_output_b_valid           (io_output_b_valid                         ), //i
    .io_output_b_ready           (writeOnly_io_output_b_ready               ), //o
    .io_output_b_payload_id      (io_output_b_payload_id[3:0]               ), //i
    .io_output_b_payload_resp    (io_output_b_payload_resp[1:0]             ), //i
    .io_axiClk                   (io_axiClk                                 ), //i
    .resetCtrl_axiReset          (resetCtrl_axiReset                        )  //i
  );
  assign io_input_ar_ready = readOnly_io_input_ar_ready;
  assign io_input_r_valid = readOnly_io_input_r_valid;
  assign io_input_r_payload_data = readOnly_io_input_r_payload_data;
  assign io_input_r_payload_id = readOnly_io_input_r_payload_id;
  assign io_input_r_payload_resp = readOnly_io_input_r_payload_resp;
  assign io_input_r_payload_last = readOnly_io_input_r_payload_last;
  assign io_input_aw_ready = writeOnly_io_input_aw_ready;
  assign io_input_w_ready = writeOnly_io_input_w_ready;
  assign io_input_b_valid = writeOnly_io_input_b_valid;
  assign io_input_b_payload_id = writeOnly_io_input_b_payload_id;
  assign io_input_b_payload_resp = writeOnly_io_input_b_payload_resp;
  assign io_output_ar_valid = readOnly_io_output_ar_valid;
  assign io_output_ar_payload_addr = readOnly_io_output_ar_payload_addr;
  assign io_output_ar_payload_id = readOnly_io_output_ar_payload_id;
  assign io_output_ar_payload_region = readOnly_io_output_ar_payload_region;
  assign io_output_ar_payload_len = readOnly_io_output_ar_payload_len;
  assign io_output_ar_payload_size = readOnly_io_output_ar_payload_size;
  assign io_output_ar_payload_burst = readOnly_io_output_ar_payload_burst;
  assign io_output_ar_payload_lock = readOnly_io_output_ar_payload_lock;
  assign io_output_ar_payload_cache = readOnly_io_output_ar_payload_cache;
  assign io_output_ar_payload_qos = readOnly_io_output_ar_payload_qos;
  assign io_output_ar_payload_prot = readOnly_io_output_ar_payload_prot;
  assign io_output_r_ready = readOnly_io_output_r_ready;
  assign io_output_aw_valid = writeOnly_io_output_aw_valid;
  assign io_output_aw_payload_addr = writeOnly_io_output_aw_payload_addr;
  assign io_output_aw_payload_id = writeOnly_io_output_aw_payload_id;
  assign io_output_aw_payload_region = writeOnly_io_output_aw_payload_region;
  assign io_output_aw_payload_len = writeOnly_io_output_aw_payload_len;
  assign io_output_aw_payload_size = writeOnly_io_output_aw_payload_size;
  assign io_output_aw_payload_burst = writeOnly_io_output_aw_payload_burst;
  assign io_output_aw_payload_lock = writeOnly_io_output_aw_payload_lock;
  assign io_output_aw_payload_cache = writeOnly_io_output_aw_payload_cache;
  assign io_output_aw_payload_qos = writeOnly_io_output_aw_payload_qos;
  assign io_output_aw_payload_prot = writeOnly_io_output_aw_payload_prot;
  assign io_output_w_valid = writeOnly_io_output_w_valid;
  assign io_output_w_payload_data = writeOnly_io_output_w_payload_data;
  assign io_output_w_payload_strb = writeOnly_io_output_w_payload_strb;
  assign io_output_w_payload_last = writeOnly_io_output_w_payload_last;
  assign io_output_b_ready = writeOnly_io_output_b_ready;

endmodule

module DandRiscvSimple (
  output reg          icache_ar_valid,
  input               icache_ar_ready,
  output reg [63:0]   icache_ar_payload_addr,
  output reg [1:0]    icache_ar_payload_id,
  output reg [7:0]    icache_ar_payload_len,
  output reg [2:0]    icache_ar_payload_size,
  output reg [1:0]    icache_ar_payload_burst,
  input               icache_r_valid,
  output              icache_r_ready,
  input      [63:0]   icache_r_payload_data,
  input      [1:0]    icache_r_payload_id,
  input      [1:0]    icache_r_payload_resp,
  input               icache_r_payload_last,
  output reg          dcache_ar_valid,
  input               dcache_ar_ready,
  output reg [63:0]   dcache_ar_payload_addr,
  output reg [1:0]    dcache_ar_payload_id,
  output reg [7:0]    dcache_ar_payload_len,
  output reg [2:0]    dcache_ar_payload_size,
  output reg [1:0]    dcache_ar_payload_burst,
  input               dcache_r_valid,
  output              dcache_r_ready,
  input      [63:0]   dcache_r_payload_data,
  input      [1:0]    dcache_r_payload_id,
  input      [1:0]    dcache_r_payload_resp,
  input               dcache_r_payload_last,
  output reg          dcache_aw_valid,
  input               dcache_aw_ready,
  output reg [63:0]   dcache_aw_payload_addr,
  output reg [1:0]    dcache_aw_payload_id,
  output reg [7:0]    dcache_aw_payload_len,
  output reg [2:0]    dcache_aw_payload_size,
  output reg [1:0]    dcache_aw_payload_burst,
  output reg          dcache_w_valid,
  input               dcache_w_ready,
  output reg [63:0]   dcache_w_payload_data,
  output reg [7:0]    dcache_w_payload_strb,
  output reg          dcache_w_payload_last,
  input               dcache_b_valid,
  output              dcache_b_ready,
  input      [1:0]    dcache_b_payload_id,
  input      [1:0]    dcache_b_payload_resp,
  input               io_axiClk,
  input               resetCtrl_axiReset
);
  localparam CsrCtrlEnum_IDLE = 4'd0;
  localparam CsrCtrlEnum_ECALL = 4'd1;
  localparam CsrCtrlEnum_EBREAK = 4'd2;
  localparam CsrCtrlEnum_MRET = 4'd3;
  localparam CsrCtrlEnum_CSRRW = 4'd4;
  localparam CsrCtrlEnum_CSRRS = 4'd5;
  localparam CsrCtrlEnum_CSRRC = 4'd6;
  localparam CsrCtrlEnum_CSRRWI = 4'd7;
  localparam CsrCtrlEnum_CSRRSI = 4'd8;
  localparam CsrCtrlEnum_CSRRCI = 4'd9;
  localparam AluCtrlEnum_IDLE = 5'd0;
  localparam AluCtrlEnum_ADD = 5'd1;
  localparam AluCtrlEnum_SUB = 5'd2;
  localparam AluCtrlEnum_SLT = 5'd3;
  localparam AluCtrlEnum_SLTU = 5'd4;
  localparam AluCtrlEnum_XOR_1 = 5'd5;
  localparam AluCtrlEnum_SLL_1 = 5'd6;
  localparam AluCtrlEnum_SRL_1 = 5'd7;
  localparam AluCtrlEnum_SRA_1 = 5'd8;
  localparam AluCtrlEnum_AND_1 = 5'd9;
  localparam AluCtrlEnum_OR_1 = 5'd10;
  localparam AluCtrlEnum_LUI = 5'd11;
  localparam AluCtrlEnum_AUIPC = 5'd12;
  localparam AluCtrlEnum_JAL = 5'd13;
  localparam AluCtrlEnum_JALR = 5'd14;
  localparam AluCtrlEnum_BEQ = 5'd15;
  localparam AluCtrlEnum_BNE = 5'd16;
  localparam AluCtrlEnum_BLT = 5'd17;
  localparam AluCtrlEnum_BGE = 5'd18;
  localparam AluCtrlEnum_BLTU = 5'd19;
  localparam AluCtrlEnum_BGEU = 5'd20;
  localparam AluCtrlEnum_CSR = 5'd21;
  localparam MemCtrlEnum_IDLE = 4'd0;
  localparam MemCtrlEnum_LB = 4'd1;
  localparam MemCtrlEnum_LBU = 4'd2;
  localparam MemCtrlEnum_LH = 4'd3;
  localparam MemCtrlEnum_LHU = 4'd4;
  localparam MemCtrlEnum_LW = 4'd5;
  localparam MemCtrlEnum_LWU = 4'd6;
  localparam MemCtrlEnum_LD = 4'd7;
  localparam MemCtrlEnum_SB = 4'd8;
  localparam MemCtrlEnum_SH = 4'd9;
  localparam MemCtrlEnum_SW = 4'd10;
  localparam MemCtrlEnum_SD = 4'd11;

  wire                regFileModule_1_write_ports_rd_wen;
  wire                clint_1_ecall;
  wire                clint_1_ebreak;
  wire                clint_1_mret;
  wire       [63:0]   timer_1_addr;
  wire                iCache_1_next_level_rsp_valid;
  wire                dCache_1_next_level_rsp_valid;
  wire                dCache_1_next_level_rsp_payload_rvalid;
  wire                dCache_1_cpu_bypass_rsp_valid;
  wire                fetch_FetchPlugin_pc_stream_fifo_ports_m_ports_valid;
  wire       [63:0]   fetch_FetchPlugin_pc_stream_fifo_ports_m_ports_payload;
  wire                fetch_FetchPlugin_pc_stream_fifo_ports_s_ports_ready;
  wire       [63:0]   fetch_FetchPlugin_pc_stream_fifo_next_payload;
  wire                fetch_FetchPlugin_pc_stream_fifo_next_valid;
  wire                fetch_FetchPlugin_predict_taken_fifo_ports_m_ports_valid;
  wire                fetch_FetchPlugin_predict_taken_fifo_ports_m_ports_payload;
  wire                fetch_FetchPlugin_predict_taken_fifo_ports_s_ports_ready;
  wire                fetch_FetchPlugin_instruction_stream_fifo_ports_m_ports_valid;
  wire       [31:0]   fetch_FetchPlugin_instruction_stream_fifo_ports_m_ports_payload;
  wire                fetch_FetchPlugin_instruction_stream_fifo_ports_s_ports_ready;
  wire                gshare_predictor_1_predict_taken;
  wire       [4:0]    gshare_predictor_1_predict_history;
  wire       [63:0]   gshare_predictor_1_predict_pc_next;
  wire       [63:0]   regFileModule_1_read_ports_rs1_value;
  wire       [63:0]   regFileModule_1_read_ports_rs2_value;
  wire       [63:0]   csrRegfile_1_cpu_ports_rdata;
  wire       [63:0]   csrRegfile_1_clint_ports_mtvec;
  wire       [63:0]   csrRegfile_1_clint_ports_mepc;
  wire       [63:0]   csrRegfile_1_clint_ports_mstatus;
  wire                csrRegfile_1_clint_ports_global_int_en;
  wire                csrRegfile_1_clint_ports_mtime_int_en;
  wire                csrRegfile_1_clint_ports_mtime_int_pend;
  wire                clint_1_csr_ports_mepc_wen;
  wire       [63:0]   clint_1_csr_ports_mepc_wdata;
  wire                clint_1_csr_ports_mcause_wen;
  wire       [63:0]   clint_1_csr_ports_mcause_wdata;
  wire                clint_1_csr_ports_mstatus_wen;
  wire       [63:0]   clint_1_csr_ports_mstatus_wdata;
  wire                clint_1_int_en;
  wire       [63:0]   clint_1_int_pc;
  wire                clint_1_int_hold;
  wire       [63:0]   timer_1_rdata;
  wire                timer_1_timer_int;
  wire                iCache_1_cpu_cmd_ready;
  wire                iCache_1_cpu_rsp_valid;
  wire       [31:0]   iCache_1_cpu_rsp_payload_data;
  wire                iCache_1_sram_0_ports_cmd_valid;
  wire       [3:0]    iCache_1_sram_0_ports_cmd_payload_addr;
  wire       [15:0]   iCache_1_sram_0_ports_cmd_payload_wen;
  wire       [511:0]  iCache_1_sram_0_ports_cmd_payload_wdata;
  wire       [63:0]   iCache_1_sram_0_ports_cmd_payload_wstrb;
  wire                iCache_1_sram_1_ports_cmd_valid;
  wire       [3:0]    iCache_1_sram_1_ports_cmd_payload_addr;
  wire       [15:0]   iCache_1_sram_1_ports_cmd_payload_wen;
  wire       [511:0]  iCache_1_sram_1_ports_cmd_payload_wdata;
  wire       [63:0]   iCache_1_sram_1_ports_cmd_payload_wstrb;
  wire                iCache_1_sram_2_ports_cmd_valid;
  wire       [3:0]    iCache_1_sram_2_ports_cmd_payload_addr;
  wire       [15:0]   iCache_1_sram_2_ports_cmd_payload_wen;
  wire       [511:0]  iCache_1_sram_2_ports_cmd_payload_wdata;
  wire       [63:0]   iCache_1_sram_2_ports_cmd_payload_wstrb;
  wire                iCache_1_sram_3_ports_cmd_valid;
  wire       [3:0]    iCache_1_sram_3_ports_cmd_payload_addr;
  wire       [15:0]   iCache_1_sram_3_ports_cmd_payload_wen;
  wire       [511:0]  iCache_1_sram_3_ports_cmd_payload_wdata;
  wire       [63:0]   iCache_1_sram_3_ports_cmd_payload_wstrb;
  wire                iCache_1_next_level_cmd_valid;
  wire       [63:0]   iCache_1_next_level_cmd_payload_addr;
  wire       [3:0]    iCache_1_next_level_cmd_payload_len;
  wire       [2:0]    iCache_1_next_level_cmd_payload_size;
  wire                sramBanks_2_sram_0_ports_rsp_valid;
  wire       [511:0]  sramBanks_2_sram_0_ports_rsp_payload_data;
  wire                sramBanks_2_sram_1_ports_rsp_valid;
  wire       [511:0]  sramBanks_2_sram_1_ports_rsp_payload_data;
  wire                sramBanks_2_sram_2_ports_rsp_valid;
  wire       [511:0]  sramBanks_2_sram_2_ports_rsp_payload_data;
  wire                sramBanks_2_sram_3_ports_rsp_valid;
  wire       [511:0]  sramBanks_2_sram_3_ports_rsp_payload_data;
  wire                dCache_1_stall;
  wire                dCache_1_cpu_cmd_ready;
  wire                dCache_1_cpu_rsp_valid;
  wire       [63:0]   dCache_1_cpu_rsp_payload_data;
  wire                dCache_1_sram_0_ports_cmd_valid;
  wire       [1:0]    dCache_1_sram_0_ports_cmd_payload_addr;
  wire       [7:0]    dCache_1_sram_0_ports_cmd_payload_wen;
  wire       [511:0]  dCache_1_sram_0_ports_cmd_payload_wdata;
  wire       [63:0]   dCache_1_sram_0_ports_cmd_payload_wstrb;
  wire                dCache_1_sram_1_ports_cmd_valid;
  wire       [1:0]    dCache_1_sram_1_ports_cmd_payload_addr;
  wire       [7:0]    dCache_1_sram_1_ports_cmd_payload_wen;
  wire       [511:0]  dCache_1_sram_1_ports_cmd_payload_wdata;
  wire       [63:0]   dCache_1_sram_1_ports_cmd_payload_wstrb;
  wire                dCache_1_sram_2_ports_cmd_valid;
  wire       [1:0]    dCache_1_sram_2_ports_cmd_payload_addr;
  wire       [7:0]    dCache_1_sram_2_ports_cmd_payload_wen;
  wire       [511:0]  dCache_1_sram_2_ports_cmd_payload_wdata;
  wire       [63:0]   dCache_1_sram_2_ports_cmd_payload_wstrb;
  wire                dCache_1_sram_3_ports_cmd_valid;
  wire       [1:0]    dCache_1_sram_3_ports_cmd_payload_addr;
  wire       [7:0]    dCache_1_sram_3_ports_cmd_payload_wen;
  wire       [511:0]  dCache_1_sram_3_ports_cmd_payload_wdata;
  wire       [63:0]   dCache_1_sram_3_ports_cmd_payload_wstrb;
  wire                dCache_1_next_level_cmd_valid;
  wire       [63:0]   dCache_1_next_level_cmd_payload_addr;
  wire       [3:0]    dCache_1_next_level_cmd_payload_len;
  wire       [2:0]    dCache_1_next_level_cmd_payload_size;
  wire                dCache_1_next_level_cmd_payload_wen;
  wire       [63:0]   dCache_1_next_level_cmd_payload_wdata;
  wire       [7:0]    dCache_1_next_level_cmd_payload_wstrb;
  wire                dCache_1_cpu_bypass_cmd_valid;
  wire       [63:0]   dCache_1_cpu_bypass_cmd_payload_addr;
  wire                dCache_1_cpu_bypass_cmd_payload_wen;
  wire       [63:0]   dCache_1_cpu_bypass_cmd_payload_wdata;
  wire       [7:0]    dCache_1_cpu_bypass_cmd_payload_wstrb;
  wire       [2:0]    dCache_1_cpu_bypass_cmd_payload_size;
  wire                sramBanks_3_sram_0_ports_rsp_valid;
  wire       [511:0]  sramBanks_3_sram_0_ports_rsp_payload_data;
  wire                sramBanks_3_sram_1_ports_rsp_valid;
  wire       [511:0]  sramBanks_3_sram_1_ports_rsp_payload_data;
  wire                sramBanks_3_sram_2_ports_rsp_valid;
  wire       [511:0]  sramBanks_3_sram_2_ports_rsp_payload_data;
  wire                sramBanks_3_sram_3_ports_rsp_valid;
  wire       [511:0]  sramBanks_3_sram_3_ports_rsp_payload_data;
  wire       [11:0]   _zz__zz_decode_DecodePlugin_imm_2;
  wire       [11:0]   _zz__zz_decode_DecodePlugin_imm_4;
  wire       [19:0]   _zz__zz_decode_DecodePlugin_imm_6;
  wire       [31:0]   _zz__zz_decode_DecodePlugin_imm_8;
  wire       [63:0]   _zz_execute_ALUPlugin_add_result;
  wire       [63:0]   _zz_execute_ALUPlugin_add_result_1;
  wire       [63:0]   _zz_execute_ALUPlugin_sub_result;
  wire       [63:0]   _zz_execute_ALUPlugin_sub_result_1;
  wire       [63:0]   _zz_execute_ALUPlugin_slt_result;
  wire       [63:0]   _zz_execute_ALUPlugin_slt_result_1;
  wire       [63:0]   _zz_execute_ALUPlugin_sra_result;
  wire       [31:0]   _zz_execute_ALUPlugin_addw_result_2;
  wire       [31:0]   _zz_execute_ALUPlugin_subw_result_2;
  wire       [31:0]   _zz_execute_ALUPlugin_sraw_temp;
  wire       [63:0]   _zz_execute_ALUPlugin_blt_result;
  wire       [63:0]   _zz_execute_ALUPlugin_blt_result_1;
  wire       [63:0]   _zz_execute_ALUPlugin_bge_result;
  wire       [63:0]   _zz_execute_ALUPlugin_bge_result_1;
  wire       [63:0]   _zz_execute_ALUPlugin_pc_next;
  wire       [63:0]   _zz_execute_ALUPlugin_pc_next_1;
  wire       [63:0]   _zz_execute_ALUPlugin_pc_next_2;
  wire       [63:0]   _zz_execute_ALUPlugin_pc_next_3;
  wire       [63:0]   _zz_execute_ALUPlugin_pc_next_4;
  wire       [63:0]   _zz_execute_ALUPlugin_pc_next_5;
  wire       [63:0]   _zz_execute_ALUPlugin_pc_next_6;
  wire       [63:0]   _zz_execute_ALUPlugin_pc_next_7;
  wire       [63:0]   _zz_execute_ALUPlugin_pc_next_8;
  wire       [5:0]    _zz_memaccess_LSUPlugin_dcache_rdata;
  wire       [5:0]    _zz_memaccess_LSUPlugin_lsu_wdata;
  wire       [63:0]   writeback_RD;
  wire                memaccess_LSU_HOLD;
  wire                memaccess_TIMER_CEN;
  wire       [63:0]   memaccess_LSU_WDATA;
  wire                execute_INT_HOLD;
  wire       [63:0]   execute_REDIRECT_PC_NEXT;
  wire                execute_REDIRECT_VALID;
  wire                execute_IS_RET;
  wire                execute_IS_CALL;
  wire                execute_IS_JMP;
  wire       [4:0]    execute_BRANCH_HISTORY;
  wire                execute_BRANCH_TAKEN;
  wire                execute_BRANCH_OR_JUMP;
  wire                execute_BRANCH_OR_JALR;
  wire       [63:0]   execute_MEM_WDATA;
  wire       [63:0]   execute_ALU_RESULT;
  wire       [63:0]   decode_CSR_RDATA;
  wire                execute_CSR_WEN;
  wire                decode_CSR_WEN;
  wire       [11:0]   execute_CSR_ADDR;
  wire       [11:0]   decode_CSR_ADDR;
  wire       [3:0]    decode_CSR_CTRL;
  wire                execute_IS_STORE;
  wire                decode_IS_STORE;
  wire                execute_IS_LOAD;
  wire                decode_IS_LOAD;
  wire       [4:0]    writeback_RD_ADDR;
  wire       [4:0]    memaccess_RD_ADDR;
  wire       [4:0]    decode_RD_ADDR;
  wire                writeback_RD_WEN;
  wire                memaccess_RD_WEN;
  wire                execute_RD_WEN;
  wire                decode_RD_WEN;
  wire       [3:0]    execute_MEM_CTRL;
  wire       [3:0]    decode_MEM_CTRL;
  wire                decode_SRC2_IS_IMM;
  wire                decode_ALU_WORD;
  wire       [4:0]    decode_ALU_CTRL;
  wire       [4:0]    execute_RS2_ADDR;
  wire       [4:0]    decode_RS2_ADDR;
  wire       [4:0]    decode_RS1_ADDR;
  wire       [63:0]   decode_RS2;
  wire       [63:0]   decode_RS1;
  wire       [63:0]   decode_IMM;
  wire       [63:0]   fetch_INT_PC;
  wire                fetch_INT_EN;
  wire       [63:0]   fetch_PREDICT_PC;
  wire                decode_PREDICT_TAKEN;
  wire                fetch_PREDICT_TAKEN;
  wire                fetch_PREDICT_VALID;
  wire       [31:0]   memaccess_INSTRUCTION;
  wire       [31:0]   execute_INSTRUCTION;
  wire       [31:0]   fetch_INSTRUCTION;
  wire       [63:0]   decode_PC_NEXT;
  wire       [63:0]   fetch_PC_NEXT;
  wire       [63:0]   memaccess_PC;
  wire       [63:0]   fetch_PC;
  wire       [31:0]   writeback_INSTRUCTION;
  wire       [63:0]   writeback_PC;
  wire       [63:0]   writeback_ALU_RESULT;
  wire       [63:0]   writeback_LSU_RDATA;
  wire                writeback_IS_LOAD;
  wire       [3:0]    memaccess_MEM_CTRL;
  wire       [63:0]   memaccess_MEM_WDATA;
  wire                memaccess_IS_STORE;
  wire                memaccess_IS_LOAD;
  wire       [3:0]    execute_CSR_CTRL;
  wire       [63:0]   execute_SRC1;
  wire       [3:0]    _zz_ecall;
  wire       [11:0]   _zz_decode_to_execute_CSR_ADDR;
  wire                _zz_memaccess_arbitration_haltItself;
  wire                _zz_DecodePlugin_hazard_ctrl_rs1_from_mem;
  wire       [4:0]    _zz_DecodePlugin_hazard_rs2_from_mem;
  wire                _zz_DecodePlugin_hazard_rs1_from_mem;
  wire       [4:0]    _zz_DecodePlugin_hazard_rs1_from_mem_1;
  wire       [4:0]    _zz_DecodePlugin_hazard_rs1_from_mem_2;
  wire                _zz_DecodePlugin_hazard_rs1_from_mem_3;
  wire       [63:0]   execute_PC_NEXT;
  wire                execute_PREDICT_TAKEN;
  wire       [63:0]   execute_CSR_RDATA;
  wire                execute_ALU_WORD;
  wire                execute_CTRL_RS2_FROM_WB;
  wire                execute_CTRL_RS2_FROM_LOAD;
  wire                execute_CTRL_RS2_FROM_MEM;
  wire                execute_CTRL_RS1_FROM_WB;
  wire       [63:0]   _zz_execute_MEM_WDATA;
  wire                execute_CTRL_RS1_FROM_LOAD;
  wire       [63:0]   _zz_execute_MEM_WDATA_1;
  wire                execute_CTRL_RS1_FROM_MEM;
  wire       [63:0]   execute_RS2;
  wire                execute_RS2_FROM_WB;
  wire                execute_RS2_FROM_LOAD;
  wire                execute_RS2_FROM_MEM;
  wire       [63:0]   execute_IMM;
  wire                execute_SRC2_IS_IMM;
  wire       [63:0]   execute_RS1;
  wire                execute_RS1_FROM_WB;
  wire       [63:0]   memaccess_LSU_RDATA;
  wire                execute_RS1_FROM_LOAD;
  wire       [63:0]   memaccess_ALU_RESULT;
  wire                execute_RS1_FROM_MEM;
  wire       [63:0]   execute_PC;
  wire       [4:0]    execute_RS1_ADDR;
  wire       [4:0]    execute_RD_ADDR;
  wire       [4:0]    execute_ALU_CTRL;
  wire       [63:0]   _zz_execute_MEM_WDATA_2;
  wire       [4:0]    _zz_DecodePlugin_hazard_rs1_from_wb;
  wire                _zz_DecodePlugin_hazard_rs1_from_wb_1;
  wire       [31:0]   decode_INSTRUCTION;
  wire       [63:0]   decode_PC;
  wire       [63:0]   _zz_execute_to_memaccess_PC;
  wire       [63:0]   fetch_BPU_PC_NEXT;
  wire       [63:0]   _zz_pc_next;
  wire                when_FetchPlugin_l97;
  wire                fetch_BPU_BRANCH_TAKEN;
  wire                when_FetchPlugin_l94;
  wire                fetch_arbitration_haltItself;
  wire                fetch_arbitration_haltByOther;
  reg                 fetch_arbitration_removeIt;
  wire                fetch_arbitration_flushIt;
  wire                fetch_arbitration_flushNext;
  wire                fetch_arbitration_isValid;
  wire                fetch_arbitration_isStuck;
  wire                fetch_arbitration_isStuckByOthers;
  wire                fetch_arbitration_isFlushed;
  wire                fetch_arbitration_isMoving;
  wire                fetch_arbitration_isFiring;
  wire                decode_arbitration_haltItself;
  wire                decode_arbitration_haltByOther;
  reg                 decode_arbitration_removeIt;
  wire                decode_arbitration_flushIt;
  wire                decode_arbitration_flushNext;
  reg                 decode_arbitration_isValid;
  wire                decode_arbitration_isStuck;
  wire                decode_arbitration_isStuckByOthers;
  wire                decode_arbitration_isFlushed;
  wire                decode_arbitration_isMoving;
  wire                decode_arbitration_isFiring;
  wire                execute_arbitration_haltItself;
  wire                execute_arbitration_haltByOther;
  reg                 execute_arbitration_removeIt;
  wire                execute_arbitration_flushIt;
  wire                execute_arbitration_flushNext;
  reg                 execute_arbitration_isValid;
  wire                execute_arbitration_isStuck;
  wire                execute_arbitration_isStuckByOthers;
  wire                execute_arbitration_isFlushed;
  wire                execute_arbitration_isMoving;
  wire                execute_arbitration_isFiring;
  wire                memaccess_arbitration_haltItself;
  wire                memaccess_arbitration_haltByOther;
  reg                 memaccess_arbitration_removeIt;
  wire                memaccess_arbitration_flushIt;
  wire                memaccess_arbitration_flushNext;
  reg                 memaccess_arbitration_isValid;
  wire                memaccess_arbitration_isStuck;
  wire                memaccess_arbitration_isStuckByOthers;
  wire                memaccess_arbitration_isFlushed;
  wire                memaccess_arbitration_isMoving;
  wire                memaccess_arbitration_isFiring;
  wire                writeback_arbitration_haltItself;
  wire                writeback_arbitration_haltByOther;
  reg                 writeback_arbitration_removeIt;
  wire                writeback_arbitration_flushIt;
  wire                writeback_arbitration_flushNext;
  reg                 writeback_arbitration_isValid;
  wire                writeback_arbitration_isStuck;
  wire                writeback_arbitration_isStuckByOthers;
  wire                writeback_arbitration_isFlushed;
  wire                writeback_arbitration_isMoving;
  wire                writeback_arbitration_isFiring;
  wire                DecodePlugin_hazard_decode_rs1_req;
  wire                DecodePlugin_hazard_decode_rs2_req;
  wire       [4:0]    DecodePlugin_hazard_decode_rs1_addr;
  wire       [4:0]    DecodePlugin_hazard_decode_rs2_addr;
  wire                DecodePlugin_hazard_rs1_from_mem;
  wire                DecodePlugin_hazard_rs2_from_mem;
  wire                DecodePlugin_hazard_rs1_from_load;
  wire                DecodePlugin_hazard_rs2_from_load;
  wire                DecodePlugin_hazard_rs1_from_wb;
  wire                DecodePlugin_hazard_rs2_from_wb;
  wire                DecodePlugin_hazard_load_use;
  wire                DecodePlugin_hazard_ctrl_rs1_from_mem;
  wire                DecodePlugin_hazard_ctrl_rs2_from_mem;
  wire                DecodePlugin_hazard_ctrl_rs1_from_load;
  wire                DecodePlugin_hazard_ctrl_rs2_from_load;
  wire                DecodePlugin_hazard_ctrl_rs1_from_wb;
  wire                DecodePlugin_hazard_ctrl_rs2_from_wb;
  wire                DecodePlugin_hazard_ctrl_load_use;
  wire                ICachePlugin_icache_access_cmd_valid;
  wire                ICachePlugin_icache_access_cmd_ready;
  wire       [63:0]   ICachePlugin_icache_access_cmd_payload_addr;
  wire                ICachePlugin_icache_access_rsp_valid;
  wire       [31:0]   ICachePlugin_icache_access_rsp_payload_data;
  wire                DCachePlugin_dcache_access_cmd_valid;
  wire                DCachePlugin_dcache_access_cmd_ready;
  wire       [63:0]   DCachePlugin_dcache_access_cmd_payload_addr;
  wire                DCachePlugin_dcache_access_cmd_payload_wen;
  wire       [63:0]   DCachePlugin_dcache_access_cmd_payload_wdata;
  wire       [7:0]    DCachePlugin_dcache_access_cmd_payload_wstrb;
  wire       [2:0]    DCachePlugin_dcache_access_cmd_payload_size;
  wire                DCachePlugin_dcache_access_rsp_valid;
  wire       [63:0]   DCachePlugin_dcache_access_rsp_payload_data;
  wire                DCachePlugin_dcache_access_stall;
  reg        [63:0]   pc_next;
  reg                 fetch_valid;
  reg                 rsp_flush;
  wire                fetch_FetchPlugin_fetch_flush;
  wire                ICachePlugin_icache_access_cmd_fire;
  wire                fetch_FetchPlugin_bpu_predict_taken;
  wire                fetch_FetchPlugin_pc_in_stream_valid;
  wire                fetch_FetchPlugin_pc_in_stream_ready;
  wire       [63:0]   fetch_FetchPlugin_pc_in_stream_payload;
  wire                fetch_FetchPlugin_pc_out_stream_valid;
  wire                fetch_FetchPlugin_pc_out_stream_ready;
  wire       [63:0]   fetch_FetchPlugin_pc_out_stream_payload;
  wire                fetch_FetchPlugin_predict_taken_in_valid;
  wire                fetch_FetchPlugin_predict_taken_in_ready;
  wire                fetch_FetchPlugin_predict_taken_in_payload;
  wire                fetch_FetchPlugin_predict_taken_out_valid;
  wire                fetch_FetchPlugin_predict_taken_out_ready;
  wire                fetch_FetchPlugin_predict_taken_out_payload;
  wire                fetch_FetchPlugin_instruction_in_stream_valid;
  wire                fetch_FetchPlugin_instruction_in_stream_ready;
  wire       [31:0]   fetch_FetchPlugin_instruction_in_stream_payload;
  wire                fetch_FetchPlugin_instruction_out_stream_valid;
  wire                fetch_FetchPlugin_instruction_out_stream_ready;
  wire       [31:0]   fetch_FetchPlugin_instruction_out_stream_payload;
  wire                fetch_FetchPlugin_fifo_all_valid;
  wire       [1:0]    IDLE;
  wire       [1:0]    FETCH;
  wire       [1:0]    HALT;
  reg        [1:0]    fetch_state_next;
  reg        [1:0]    fetch_state;
  wire                when_FetchPlugin_l64;
  wire                ICachePlugin_icache_access_cmd_isStall;
  wire                when_FetchPlugin_l72;
  wire                when_FetchPlugin_l80;
  wire                when_FetchPlugin_l93;
  wire                when_FetchPlugin_l109;
  wire                ICachePlugin_icache_access_cmd_fire_1;
  wire                ICachePlugin_icache_access_cmd_fire_2;
  wire                ICachePlugin_icache_access_cmd_fire_3;
  wire                ICachePlugin_icache_access_cmd_fire_4;
  reg        [63:0]   decode_DecodePlugin_imm;
  wire       [63:0]   decode_DecodePlugin_rs1;
  wire       [63:0]   decode_DecodePlugin_rs2;
  wire                decode_DecodePlugin_rs1_req;
  wire                decode_DecodePlugin_rs2_req;
  wire       [4:0]    decode_DecodePlugin_rs1_addr;
  wire       [4:0]    decode_DecodePlugin_rs2_addr;
  wire                decode_DecodePlugin_rd_wen;
  wire       [4:0]    decode_DecodePlugin_rd_addr;
  reg        [4:0]    decode_DecodePlugin_alu_ctrl;
  wire                decode_DecodePlugin_alu_word;
  wire                decode_DecodePlugin_src2_is_imm;
  reg        [3:0]    decode_DecodePlugin_mem_ctrl;
  reg                 decode_DecodePlugin_is_load;
  reg                 decode_DecodePlugin_is_store;
  reg        [3:0]    decode_DecodePlugin_csr_ctrl;
  wire       [11:0]   decode_DecodePlugin_csr_addr;
  wire                decode_DecodePlugin_csr_wen;
  wire                when_DecodePlugin_l116;
  wire                _zz_decode_DecodePlugin_imm;
  reg        [51:0]   _zz_decode_DecodePlugin_imm_1;
  wire                _zz_decode_DecodePlugin_imm_2;
  reg        [51:0]   _zz_decode_DecodePlugin_imm_3;
  wire                _zz_decode_DecodePlugin_imm_4;
  reg        [50:0]   _zz_decode_DecodePlugin_imm_5;
  wire                _zz_decode_DecodePlugin_imm_6;
  reg        [42:0]   _zz_decode_DecodePlugin_imm_7;
  wire                _zz_decode_DecodePlugin_imm_8;
  reg        [31:0]   _zz_decode_DecodePlugin_imm_9;
  wire                _zz_decode_DecodePlugin_imm_10;
  reg        [51:0]   _zz_decode_DecodePlugin_imm_11;
  wire                when_DecodePlugin_l119;
  wire                when_DecodePlugin_l122;
  wire                when_DecodePlugin_l125;
  wire                when_DecodePlugin_l128;
  reg        [63:0]   execute_ALUPlugin_src1;
  reg        [63:0]   execute_ALUPlugin_src2;
  wire       [31:0]   execute_ALUPlugin_src1_word;
  wire       [31:0]   execute_ALUPlugin_src2_word;
  wire       [5:0]    execute_ALUPlugin_shift_bits;
  wire       [63:0]   execute_ALUPlugin_add_result;
  wire       [63:0]   execute_ALUPlugin_sub_result;
  wire                execute_ALUPlugin_slt_result;
  wire                execute_ALUPlugin_sltu_result;
  wire       [63:0]   execute_ALUPlugin_xor_result;
  wire       [63:0]   execute_ALUPlugin_sll_result;
  wire       [63:0]   execute_ALUPlugin_srl_result;
  wire       [63:0]   execute_ALUPlugin_sra_result;
  wire       [63:0]   execute_ALUPlugin_and_result;
  wire       [63:0]   execute_ALUPlugin_or_result;
  wire                _zz_execute_ALUPlugin_addw_result;
  reg        [31:0]   _zz_execute_ALUPlugin_addw_result_1;
  wire       [63:0]   execute_ALUPlugin_addw_result;
  wire                _zz_execute_ALUPlugin_subw_result;
  reg        [31:0]   _zz_execute_ALUPlugin_subw_result_1;
  wire       [63:0]   execute_ALUPlugin_subw_result;
  wire       [31:0]   execute_ALUPlugin_sllw_temp;
  wire                _zz_execute_ALUPlugin_sllw_result;
  reg        [31:0]   _zz_execute_ALUPlugin_sllw_result_1;
  wire       [63:0]   execute_ALUPlugin_sllw_result;
  wire       [31:0]   execute_ALUPlugin_srlw_temp;
  wire                _zz_execute_ALUPlugin_srlw_result;
  reg        [31:0]   _zz_execute_ALUPlugin_srlw_result_1;
  wire       [63:0]   execute_ALUPlugin_srlw_result;
  wire       [31:0]   execute_ALUPlugin_sraw_temp;
  wire                _zz_execute_ALUPlugin_sraw_result;
  reg        [31:0]   _zz_execute_ALUPlugin_sraw_result_1;
  wire       [63:0]   execute_ALUPlugin_sraw_result;
  reg        [63:0]   execute_ALUPlugin_alu_result;
  reg        [63:0]   execute_ALUPlugin_pc_next;
  wire                execute_ALUPlugin_jal;
  wire                execute_ALUPlugin_jalr;
  wire                execute_ALUPlugin_beq;
  wire                execute_ALUPlugin_bne;
  wire                execute_ALUPlugin_blt;
  wire                execute_ALUPlugin_bge;
  wire                execute_ALUPlugin_bltu;
  wire                execute_ALUPlugin_bgeu;
  wire                execute_ALUPlugin_branch_or_jalr;
  wire                execute_ALUPlugin_branch_or_jump;
  reg        [63:0]   execute_ALUPlugin_branch_src1;
  reg        [63:0]   execute_ALUPlugin_branch_src2;
  wire                execute_ALUPlugin_rd_is_link;
  wire                execute_ALUPlugin_rs1_is_link;
  reg                 execute_ALUPlugin_is_call;
  reg                 execute_ALUPlugin_is_ret;
  reg                 execute_ALUPlugin_is_jmp;
  reg        [63:0]   execute_ALUPlugin_redirect_pc_next;
  reg                 execute_ALUPlugin_redirect_valid;
  wire                when_AluPlugin_l77;
  wire                when_AluPlugin_l95;
  wire                when_AluPlugin_l146;
  wire                when_AluPlugin_l153;
  wire       [62:0]   _zz_execute_ALUPlugin_alu_result;
  wire       [62:0]   _zz_execute_ALUPlugin_alu_result_1;
  wire                when_AluPlugin_l169;
  wire                when_AluPlugin_l176;
  wire                when_AluPlugin_l183;
  wire                execute_ALUPlugin_beq_result;
  wire                execute_ALUPlugin_bne_result;
  wire                execute_ALUPlugin_blt_result;
  wire                execute_ALUPlugin_bge_result;
  wire                execute_ALUPlugin_bltu_result;
  wire                execute_ALUPlugin_bgeu_result;
  wire                execute_ALUPlugin_branch_taken;
  reg        [4:0]    execute_ALUPlugin_branch_history;
  wire                when_AluPlugin_l226;
  wire                when_AluPlugin_l234;
  wire                when_AluPlugin_l270;
  reg        [63:0]   execute_ExcepPlugin_csr_wdata;
  wire       [63:0]   execute_ExcepPlugin_csrrs_wdata;
  wire       [63:0]   execute_ExcepPlugin_csrrc_wdata;
  wire       [63:0]   execute_ExcepPlugin_csrrsi_wdata;
  wire       [63:0]   execute_ExcepPlugin_csrrci_wdata;
  wire       [63:0]   memaccess_LSUPlugin_cpu_addr;
  wire       [2:0]    memaccess_LSUPlugin_cpu_addr_offset;
  wire                memaccess_LSUPlugin_is_mem;
  wire                memaccess_LSUPlugin_is_timer;
  wire       [63:0]   memaccess_LSUPlugin_dcache_rdata;
  wire                _zz_memaccess_LSUPlugin_dcache_lb;
  reg        [55:0]   _zz_memaccess_LSUPlugin_dcache_lb_1;
  wire       [63:0]   memaccess_LSUPlugin_dcache_lb;
  reg        [55:0]   _zz_memaccess_LSUPlugin_dcache_lbu;
  wire       [63:0]   memaccess_LSUPlugin_dcache_lbu;
  wire                _zz_memaccess_LSUPlugin_dcache_lh;
  reg        [47:0]   _zz_memaccess_LSUPlugin_dcache_lh_1;
  wire       [63:0]   memaccess_LSUPlugin_dcache_lh;
  reg        [47:0]   _zz_memaccess_LSUPlugin_dcache_lhu;
  wire       [63:0]   memaccess_LSUPlugin_dcache_lhu;
  wire                _zz_memaccess_LSUPlugin_dcache_lw;
  reg        [31:0]   _zz_memaccess_LSUPlugin_dcache_lw_1;
  wire       [63:0]   memaccess_LSUPlugin_dcache_lw;
  reg        [31:0]   _zz_memaccess_LSUPlugin_dcache_lwu;
  wire       [63:0]   memaccess_LSUPlugin_dcache_lwu;
  reg        [63:0]   memaccess_LSUPlugin_dcache_data_load;
  wire                _zz_memaccess_LSUPlugin_dcache_sb;
  reg        [55:0]   _zz_memaccess_LSUPlugin_dcache_sb_1;
  wire       [63:0]   memaccess_LSUPlugin_dcache_sb;
  wire                _zz_memaccess_LSUPlugin_dcache_sh;
  reg        [47:0]   _zz_memaccess_LSUPlugin_dcache_sh_1;
  wire       [63:0]   memaccess_LSUPlugin_dcache_sh;
  wire                _zz_memaccess_LSUPlugin_dcache_sw;
  reg        [31:0]   _zz_memaccess_LSUPlugin_dcache_sw_1;
  wire       [63:0]   memaccess_LSUPlugin_dcache_sw;
  reg        [63:0]   memaccess_LSUPlugin_dcache_wdata;
  reg        [7:0]    memaccess_LSUPlugin_dcache_wstrb;
  wire                memaccess_LSUPlugin_lsu_ready;
  wire       [63:0]   memaccess_LSUPlugin_lsu_addr;
  wire       [63:0]   memaccess_LSUPlugin_lsu_rdata;
  wire       [63:0]   memaccess_LSUPlugin_lsu_wdata;
  wire                memaccess_LSUPlugin_lsu_wen;
  wire       [7:0]    memaccess_LSUPlugin_lsu_wstrb;
  reg        [2:0]    memaccess_LSUPlugin_lsu_size;
  reg        [7:0]    _zz_memaccess_LSUPlugin_dcache_wstrb;
  reg        [7:0]    _zz_memaccess_LSUPlugin_dcache_wstrb_1;
  reg        [7:0]    _zz_memaccess_LSUPlugin_dcache_wstrb_2;
  wire       [7:0]    _zz_memaccess_LSUPlugin_dcache_wstrb_3;
  reg        [3:0]    ar_len_cnt;
  wire                icache_ar_fire;
  wire                when_ICachePlugin_l141;
  wire                when_ICachePlugin_l149;
  wire                icache_ar_fire_1;
  wire                icache_ar_fire_2;
  reg                 _zz_when_DCachePlugin_l349;
  reg        [3:0]    _zz_when_DCachePlugin_l258;
  wire                when_DCachePlugin_l265;
  wire                when_DCachePlugin_l313;
  wire                when_DCachePlugin_l267;
  wire                when_DCachePlugin_l233;
  reg                 _zz_cpu_bypass_rsp_valid;
  reg                 _zz_cpu_bypass_rsp_valid_1;
  wire                when_DCachePlugin_l239;
  wire                when_DCachePlugin_l254;
  wire                when_DCachePlugin_l258;
  wire                dcache_ar_fire;
  wire                dcache_ar_fire_1;
  wire                when_DCachePlugin_l269;
  wire                dcache_ar_fire_2;
  wire                when_DCachePlugin_l303;
  wire                dcache_aw_fire;
  wire                when_DCachePlugin_l335;
  wire                dcache_w_fire;
  wire                when_DCachePlugin_l349;
  wire                dcache_aw_fire_1;
  wire                dcache_w_fire_1;
  wire                when_DCachePlugin_l350;
  wire                dcache_aw_fire_2;
  wire                dcache_w_fire_2;
  wire                when_DCachePlugin_l352;
  wire                dcache_aw_fire_3;
  wire                dcache_w_fire_3;
  wire                when_DCachePlugin_l357;
  wire                when_DCachePlugin_l356;
  wire                dcache_aw_fire_4;
  wire                dcache_w_fire_4;
  wire                dcache_aw_fire_5;
  wire                dcache_w_fire_5;
  wire                when_Pipeline_l127;
  reg        [63:0]   fetch_to_decode_PC;
  wire                when_Pipeline_l127_1;
  reg        [63:0]   decode_to_execute_PC;
  wire                when_Pipeline_l127_2;
  reg        [63:0]   execute_to_memaccess_PC;
  wire                when_Pipeline_l127_3;
  reg        [63:0]   memaccess_to_writeback_PC;
  wire                when_Pipeline_l127_4;
  reg        [63:0]   fetch_to_decode_PC_NEXT;
  wire                when_Pipeline_l127_5;
  reg        [63:0]   decode_to_execute_PC_NEXT;
  wire                when_Pipeline_l127_6;
  reg        [31:0]   fetch_to_decode_INSTRUCTION;
  wire                when_Pipeline_l127_7;
  reg        [31:0]   decode_to_execute_INSTRUCTION;
  wire                when_Pipeline_l127_8;
  reg        [31:0]   execute_to_memaccess_INSTRUCTION;
  wire                when_Pipeline_l127_9;
  reg        [31:0]   memaccess_to_writeback_INSTRUCTION;
  wire                when_Pipeline_l127_10;
  reg                 fetch_to_decode_PREDICT_TAKEN;
  wire                when_Pipeline_l127_11;
  reg                 decode_to_execute_PREDICT_TAKEN;
  wire                when_Pipeline_l127_12;
  reg        [63:0]   decode_to_execute_IMM;
  wire                when_Pipeline_l127_13;
  reg        [63:0]   decode_to_execute_RS1;
  wire                when_Pipeline_l127_14;
  reg        [63:0]   decode_to_execute_RS2;
  wire                when_Pipeline_l127_15;
  reg        [4:0]    decode_to_execute_RS1_ADDR;
  wire                when_Pipeline_l127_16;
  reg        [4:0]    decode_to_execute_RS2_ADDR;
  wire                when_Pipeline_l127_17;
  reg        [4:0]    decode_to_execute_ALU_CTRL;
  wire                when_Pipeline_l127_18;
  reg                 decode_to_execute_ALU_WORD;
  wire                when_Pipeline_l127_19;
  reg                 decode_to_execute_SRC2_IS_IMM;
  wire                when_Pipeline_l127_20;
  reg        [3:0]    decode_to_execute_MEM_CTRL;
  wire                when_Pipeline_l127_21;
  reg        [3:0]    execute_to_memaccess_MEM_CTRL;
  wire                when_Pipeline_l127_22;
  reg                 decode_to_execute_RD_WEN;
  wire                when_Pipeline_l127_23;
  reg                 execute_to_memaccess_RD_WEN;
  wire                when_Pipeline_l127_24;
  reg                 memaccess_to_writeback_RD_WEN;
  wire                when_Pipeline_l127_25;
  reg        [4:0]    decode_to_execute_RD_ADDR;
  wire                when_Pipeline_l127_26;
  reg        [4:0]    execute_to_memaccess_RD_ADDR;
  wire                when_Pipeline_l127_27;
  reg        [4:0]    memaccess_to_writeback_RD_ADDR;
  wire                when_Pipeline_l127_28;
  reg                 decode_to_execute_IS_LOAD;
  wire                when_Pipeline_l127_29;
  reg                 execute_to_memaccess_IS_LOAD;
  wire                when_Pipeline_l127_30;
  reg                 memaccess_to_writeback_IS_LOAD;
  wire                when_Pipeline_l127_31;
  reg                 decode_to_execute_IS_STORE;
  wire                when_Pipeline_l127_32;
  reg                 execute_to_memaccess_IS_STORE;
  wire                when_Pipeline_l127_33;
  reg        [3:0]    decode_to_execute_CSR_CTRL;
  wire                when_Pipeline_l127_34;
  reg        [11:0]   decode_to_execute_CSR_ADDR;
  wire                when_Pipeline_l127_35;
  reg                 decode_to_execute_CSR_WEN;
  wire                when_Pipeline_l127_36;
  reg        [63:0]   decode_to_execute_CSR_RDATA;
  wire                when_Pipeline_l127_37;
  reg        [63:0]   execute_to_memaccess_ALU_RESULT;
  wire                when_Pipeline_l127_38;
  reg        [63:0]   memaccess_to_writeback_ALU_RESULT;
  wire                when_Pipeline_l127_39;
  reg        [63:0]   execute_to_memaccess_MEM_WDATA;
  wire                when_Pipeline_l127_40;
  reg        [63:0]   memaccess_to_writeback_LSU_RDATA;
  wire                when_Pipeline_l163;
  wire                when_Pipeline_l166;
  wire                when_Pipeline_l163_1;
  wire                when_Pipeline_l166_1;
  wire                when_Pipeline_l163_2;
  wire                when_Pipeline_l166_2;
  wire                when_Pipeline_l163_3;
  wire                when_Pipeline_l166_3;
  function [55:0] zz__zz_memaccess_LSUPlugin_dcache_lbu(input dummy);
    begin
      zz__zz_memaccess_LSUPlugin_dcache_lbu[55] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[54] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[53] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[52] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[51] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[50] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[49] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[48] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[47] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[46] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[45] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[44] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[43] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[42] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[41] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[40] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[39] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[38] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[37] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[36] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[35] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[34] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[33] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[32] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[31] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[30] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[29] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[28] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[27] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[26] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[25] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[24] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[23] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[22] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[21] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[20] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[19] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[18] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[17] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[16] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[15] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[14] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[13] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[12] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[11] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[10] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[9] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[8] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[7] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[6] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[5] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[4] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[3] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[2] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[1] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[0] = 1'b0;
    end
  endfunction
  wire [55:0] _zz_1;
  function [47:0] zz__zz_memaccess_LSUPlugin_dcache_lhu(input dummy);
    begin
      zz__zz_memaccess_LSUPlugin_dcache_lhu[47] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[46] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[45] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[44] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[43] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[42] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[41] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[40] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[39] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[38] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[37] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[36] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[35] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[34] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[33] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[32] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[31] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[30] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[29] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[28] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[27] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[26] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[25] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[24] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[23] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[22] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[21] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[20] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[19] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[18] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[17] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[16] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[15] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[14] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[13] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[12] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[11] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[10] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[9] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[8] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[7] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[6] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[5] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[4] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[3] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[2] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[1] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[0] = 1'b0;
    end
  endfunction
  wire [47:0] _zz_2;
  function [31:0] zz__zz_memaccess_LSUPlugin_dcache_lwu(input dummy);
    begin
      zz__zz_memaccess_LSUPlugin_dcache_lwu[31] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[30] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[29] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[28] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[27] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[26] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[25] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[24] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[23] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[22] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[21] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[20] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[19] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[18] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[17] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[16] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[15] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[14] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[13] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[12] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[11] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[10] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[9] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[8] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[7] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[6] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[5] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[4] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[3] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[2] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[1] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[0] = 1'b0;
    end
  endfunction
  wire [31:0] _zz_3;
  function [7:0] zz__zz_memaccess_LSUPlugin_dcache_wstrb(input dummy);
    begin
      zz__zz_memaccess_LSUPlugin_dcache_wstrb = 8'h0;
      zz__zz_memaccess_LSUPlugin_dcache_wstrb[0] = 1'b1;
    end
  endfunction
  wire [7:0] _zz_4;
  function [7:0] zz__zz_memaccess_LSUPlugin_dcache_wstrb_1(input dummy);
    begin
      zz__zz_memaccess_LSUPlugin_dcache_wstrb_1 = 8'h0;
      zz__zz_memaccess_LSUPlugin_dcache_wstrb_1[1 : 0] = 2'b11;
    end
  endfunction
  wire [7:0] _zz_5;
  function [7:0] zz__zz_memaccess_LSUPlugin_dcache_wstrb_2(input dummy);
    begin
      zz__zz_memaccess_LSUPlugin_dcache_wstrb_2 = 8'h0;
      zz__zz_memaccess_LSUPlugin_dcache_wstrb_2[3 : 0] = 4'b1111;
    end
  endfunction
  wire [7:0] _zz_6;

  assign _zz__zz_decode_DecodePlugin_imm_2 = {decode_INSTRUCTION[31 : 25],decode_INSTRUCTION[11 : 7]};
  assign _zz__zz_decode_DecodePlugin_imm_4 = {{{decode_INSTRUCTION[31],decode_INSTRUCTION[7]},decode_INSTRUCTION[30 : 25]},decode_INSTRUCTION[11 : 8]};
  assign _zz__zz_decode_DecodePlugin_imm_6 = {{{decode_INSTRUCTION[31],decode_INSTRUCTION[19 : 12]},decode_INSTRUCTION[20]},decode_INSTRUCTION[30 : 21]};
  assign _zz__zz_decode_DecodePlugin_imm_8 = {decode_INSTRUCTION[31 : 12],12'h0};
  assign _zz_execute_ALUPlugin_add_result = execute_ALUPlugin_src1;
  assign _zz_execute_ALUPlugin_add_result_1 = execute_ALUPlugin_src2;
  assign _zz_execute_ALUPlugin_sub_result = execute_ALUPlugin_src1;
  assign _zz_execute_ALUPlugin_sub_result_1 = execute_ALUPlugin_src2;
  assign _zz_execute_ALUPlugin_slt_result = execute_ALUPlugin_src1;
  assign _zz_execute_ALUPlugin_slt_result_1 = execute_ALUPlugin_src2;
  assign _zz_execute_ALUPlugin_sra_result = execute_ALUPlugin_src1;
  assign _zz_execute_ALUPlugin_addw_result_2 = execute_ALUPlugin_add_result[31 : 0];
  assign _zz_execute_ALUPlugin_subw_result_2 = execute_ALUPlugin_sub_result[31 : 0];
  assign _zz_execute_ALUPlugin_sraw_temp = execute_ALUPlugin_src1_word;
  assign _zz_execute_ALUPlugin_blt_result = execute_ALUPlugin_branch_src1;
  assign _zz_execute_ALUPlugin_blt_result_1 = execute_ALUPlugin_branch_src2;
  assign _zz_execute_ALUPlugin_bge_result = execute_ALUPlugin_branch_src2;
  assign _zz_execute_ALUPlugin_bge_result_1 = execute_ALUPlugin_branch_src1;
  assign _zz_execute_ALUPlugin_pc_next = (_zz_execute_ALUPlugin_pc_next_1 & _zz_execute_ALUPlugin_pc_next_4);
  assign _zz_execute_ALUPlugin_pc_next_1 = ($signed(_zz_execute_ALUPlugin_pc_next_2) + $signed(_zz_execute_ALUPlugin_pc_next_3));
  assign _zz_execute_ALUPlugin_pc_next_2 = execute_ALUPlugin_branch_src1;
  assign _zz_execute_ALUPlugin_pc_next_3 = execute_IMM;
  assign _zz_execute_ALUPlugin_pc_next_4 = (~ _zz_execute_ALUPlugin_pc_next_5);
  assign _zz_execute_ALUPlugin_pc_next_5 = 64'h0000000000000001;
  assign _zz_execute_ALUPlugin_pc_next_6 = ($signed(_zz_execute_ALUPlugin_pc_next_7) + $signed(_zz_execute_ALUPlugin_pc_next_8));
  assign _zz_execute_ALUPlugin_pc_next_7 = execute_PC;
  assign _zz_execute_ALUPlugin_pc_next_8 = execute_IMM;
  assign _zz_memaccess_LSUPlugin_dcache_rdata = ({3'd0,memaccess_LSUPlugin_cpu_addr_offset} <<< 3);
  assign _zz_memaccess_LSUPlugin_lsu_wdata = ({3'd0,memaccess_LSUPlugin_cpu_addr_offset} <<< 3);
  FIFO fetch_FetchPlugin_pc_stream_fifo (
    .ports_s_ports_valid   (fetch_FetchPlugin_pc_in_stream_valid                        ), //i
    .ports_s_ports_ready   (fetch_FetchPlugin_pc_stream_fifo_ports_s_ports_ready        ), //o
    .ports_s_ports_payload (fetch_FetchPlugin_pc_in_stream_payload[63:0]                ), //i
    .ports_m_ports_valid   (fetch_FetchPlugin_pc_stream_fifo_ports_m_ports_valid        ), //o
    .ports_m_ports_ready   (fetch_FetchPlugin_pc_out_stream_ready                       ), //i
    .ports_m_ports_payload (fetch_FetchPlugin_pc_stream_fifo_ports_m_ports_payload[63:0]), //o
    .flush                 (fetch_FetchPlugin_fetch_flush                               ), //i
    .next_payload          (fetch_FetchPlugin_pc_stream_fifo_next_payload[63:0]         ), //o
    .next_valid            (fetch_FetchPlugin_pc_stream_fifo_next_valid                 ), //o
    .io_axiClk             (io_axiClk                                                   ), //i
    .resetCtrl_axiReset    (resetCtrl_axiReset                                          )  //i
  );
  FIFO_1 fetch_FetchPlugin_predict_taken_fifo (
    .ports_s_ports_valid   (fetch_FetchPlugin_predict_taken_in_valid                  ), //i
    .ports_s_ports_ready   (fetch_FetchPlugin_predict_taken_fifo_ports_s_ports_ready  ), //o
    .ports_s_ports_payload (fetch_FetchPlugin_predict_taken_in_payload                ), //i
    .ports_m_ports_valid   (fetch_FetchPlugin_predict_taken_fifo_ports_m_ports_valid  ), //o
    .ports_m_ports_ready   (fetch_FetchPlugin_predict_taken_out_ready                 ), //i
    .ports_m_ports_payload (fetch_FetchPlugin_predict_taken_fifo_ports_m_ports_payload), //o
    .flush                 (fetch_FetchPlugin_fetch_flush                             ), //i
    .io_axiClk             (io_axiClk                                                 ), //i
    .resetCtrl_axiReset    (resetCtrl_axiReset                                        )  //i
  );
  FIFO_2 fetch_FetchPlugin_instruction_stream_fifo (
    .ports_s_ports_valid   (fetch_FetchPlugin_instruction_in_stream_valid                        ), //i
    .ports_s_ports_ready   (fetch_FetchPlugin_instruction_stream_fifo_ports_s_ports_ready        ), //o
    .ports_s_ports_payload (fetch_FetchPlugin_instruction_in_stream_payload[31:0]                ), //i
    .ports_m_ports_valid   (fetch_FetchPlugin_instruction_stream_fifo_ports_m_ports_valid        ), //o
    .ports_m_ports_ready   (fetch_FetchPlugin_instruction_out_stream_ready                       ), //i
    .ports_m_ports_payload (fetch_FetchPlugin_instruction_stream_fifo_ports_m_ports_payload[31:0]), //o
    .flush                 (fetch_FetchPlugin_fetch_flush                                        ), //i
    .io_axiClk             (io_axiClk                                                            ), //i
    .resetCtrl_axiReset    (resetCtrl_axiReset                                                   )  //i
  );
  gshare_predictor gshare_predictor_1 (
    .predict_pc         (fetch_PREDICT_PC[63:0]                  ), //i
    .predict_valid      (fetch_PREDICT_VALID                     ), //i
    .predict_taken      (gshare_predictor_1_predict_taken        ), //o
    .predict_history    (gshare_predictor_1_predict_history[4:0] ), //o
    .predict_pc_next    (gshare_predictor_1_predict_pc_next[63:0]), //o
    .train_valid        (execute_BRANCH_OR_JUMP                  ), //i
    .train_taken        (execute_BRANCH_TAKEN                    ), //i
    .train_mispredicted (when_FetchPlugin_l97                    ), //i
    .train_history      (execute_BRANCH_HISTORY[4:0]             ), //i
    .train_pc           (_zz_execute_to_memaccess_PC[63:0]       ), //i
    .train_pc_next      (_zz_pc_next[63:0]                       ), //i
    .train_is_call      (execute_IS_CALL                         ), //i
    .train_is_ret       (execute_IS_RET                          ), //i
    .train_is_jmp       (execute_IS_JMP                          ), //i
    .io_axiClk          (io_axiClk                               ), //i
    .resetCtrl_axiReset (resetCtrl_axiReset                      )  //i
  );
  RegFileModule regFileModule_1 (
    .read_ports_rs1_value (regFileModule_1_read_ports_rs1_value[63:0]), //o
    .read_ports_rs2_value (regFileModule_1_read_ports_rs2_value[63:0]), //o
    .read_ports_rs1_addr  (decode_DecodePlugin_rs1_addr[4:0]         ), //i
    .read_ports_rs2_addr  (decode_DecodePlugin_rs2_addr[4:0]         ), //i
    .read_ports_rs1_req   (decode_DecodePlugin_rs1_req               ), //i
    .read_ports_rs2_req   (decode_DecodePlugin_rs2_req               ), //i
    .write_ports_rd_value (_zz_execute_MEM_WDATA_2[63:0]             ), //i
    .write_ports_rd_addr  (_zz_DecodePlugin_hazard_rs1_from_wb[4:0]  ), //i
    .write_ports_rd_wen   (regFileModule_1_write_ports_rd_wen        ), //i
    .io_axiClk            (io_axiClk                                 ), //i
    .resetCtrl_axiReset   (resetCtrl_axiReset                        )  //i
  );
  CsrRegfile csrRegfile_1 (
    .cpu_ports_waddr            (execute_CSR_ADDR[11:0]                 ), //i
    .cpu_ports_wen              (execute_CSR_WEN                        ), //i
    .cpu_ports_wdata            (execute_ExcepPlugin_csr_wdata[63:0]    ), //i
    .cpu_ports_raddr            (_zz_decode_to_execute_CSR_ADDR[11:0]   ), //i
    .cpu_ports_rdata            (csrRegfile_1_cpu_ports_rdata[63:0]     ), //o
    .clint_ports_mepc_wen       (clint_1_csr_ports_mepc_wen             ), //i
    .clint_ports_mepc_wdata     (clint_1_csr_ports_mepc_wdata[63:0]     ), //i
    .clint_ports_mcause_wen     (clint_1_csr_ports_mcause_wen           ), //i
    .clint_ports_mcause_wdata   (clint_1_csr_ports_mcause_wdata[63:0]   ), //i
    .clint_ports_mstatus_wen    (clint_1_csr_ports_mstatus_wen          ), //i
    .clint_ports_mstatus_wdata  (clint_1_csr_ports_mstatus_wdata[63:0]  ), //i
    .clint_ports_mtvec          (csrRegfile_1_clint_ports_mtvec[63:0]   ), //o
    .clint_ports_mepc           (csrRegfile_1_clint_ports_mepc[63:0]    ), //o
    .clint_ports_mstatus        (csrRegfile_1_clint_ports_mstatus[63:0] ), //o
    .clint_ports_global_int_en  (csrRegfile_1_clint_ports_global_int_en ), //o
    .clint_ports_mtime_int_en   (csrRegfile_1_clint_ports_mtime_int_en  ), //o
    .clint_ports_mtime_int_pend (csrRegfile_1_clint_ports_mtime_int_pend), //o
    .timer_int                  (timer_1_timer_int                      ), //i
    .io_axiClk                  (io_axiClk                              ), //i
    .resetCtrl_axiReset         (resetCtrl_axiReset                     )  //i
  );
  Clint clint_1 (
    .pc                       (_zz_execute_to_memaccess_PC[63:0]      ), //i
    .pc_next                  (_zz_pc_next[63:0]                      ), //i
    .pc_next_valid            (when_FetchPlugin_l97                   ), //i
    .instruction_valid        (execute_arbitration_isValid            ), //i
    .csr_ports_mepc_wen       (clint_1_csr_ports_mepc_wen             ), //o
    .csr_ports_mepc_wdata     (clint_1_csr_ports_mepc_wdata[63:0]     ), //o
    .csr_ports_mcause_wen     (clint_1_csr_ports_mcause_wen           ), //o
    .csr_ports_mcause_wdata   (clint_1_csr_ports_mcause_wdata[63:0]   ), //o
    .csr_ports_mstatus_wen    (clint_1_csr_ports_mstatus_wen          ), //o
    .csr_ports_mstatus_wdata  (clint_1_csr_ports_mstatus_wdata[63:0]  ), //o
    .csr_ports_mtvec          (csrRegfile_1_clint_ports_mtvec[63:0]   ), //i
    .csr_ports_mepc           (csrRegfile_1_clint_ports_mepc[63:0]    ), //i
    .csr_ports_mstatus        (csrRegfile_1_clint_ports_mstatus[63:0] ), //i
    .csr_ports_global_int_en  (csrRegfile_1_clint_ports_global_int_en ), //i
    .csr_ports_mtime_int_en   (csrRegfile_1_clint_ports_mtime_int_en  ), //i
    .csr_ports_mtime_int_pend (csrRegfile_1_clint_ports_mtime_int_pend), //i
    .timer_int                (timer_1_timer_int                      ), //i
    .int_en                   (clint_1_int_en                         ), //o
    .int_pc                   (clint_1_int_pc[63:0]                   ), //o
    .int_hold                 (clint_1_int_hold                       ), //o
    .ecall                    (clint_1_ecall                          ), //i
    .ebreak                   (clint_1_ebreak                         ), //i
    .mret                     (clint_1_mret                           ), //i
    .io_axiClk                (io_axiClk                              ), //i
    .resetCtrl_axiReset       (resetCtrl_axiReset                     )  //i
  );
  Timer timer_1 (
    .cen                (memaccess_TIMER_CEN      ), //i
    .wen                (memaccess_IS_STORE       ), //i
    .addr               (timer_1_addr[63:0]       ), //i
    .wdata              (memaccess_LSU_WDATA[63:0]), //i
    .rdata              (timer_1_rdata[63:0]      ), //o
    .timer_int          (timer_1_timer_int        ), //o
    .io_axiClk          (io_axiClk                ), //i
    .resetCtrl_axiReset (resetCtrl_axiReset       )  //i
  );
  ICache iCache_1 (
    .flush                          (1'b0                                             ), //i
    .cpu_cmd_valid                  (ICachePlugin_icache_access_cmd_valid             ), //i
    .cpu_cmd_ready                  (iCache_1_cpu_cmd_ready                           ), //o
    .cpu_cmd_payload_addr           (ICachePlugin_icache_access_cmd_payload_addr[63:0]), //i
    .cpu_rsp_valid                  (iCache_1_cpu_rsp_valid                           ), //o
    .cpu_rsp_payload_data           (iCache_1_cpu_rsp_payload_data[31:0]              ), //o
    .sram_0_ports_cmd_valid         (iCache_1_sram_0_ports_cmd_valid                  ), //o
    .sram_0_ports_cmd_payload_addr  (iCache_1_sram_0_ports_cmd_payload_addr[3:0]      ), //o
    .sram_0_ports_cmd_payload_wen   (iCache_1_sram_0_ports_cmd_payload_wen[15:0]      ), //o
    .sram_0_ports_cmd_payload_wdata (iCache_1_sram_0_ports_cmd_payload_wdata[511:0]   ), //o
    .sram_0_ports_cmd_payload_wstrb (iCache_1_sram_0_ports_cmd_payload_wstrb[63:0]    ), //o
    .sram_0_ports_rsp_valid         (sramBanks_2_sram_0_ports_rsp_valid               ), //i
    .sram_0_ports_rsp_payload_data  (sramBanks_2_sram_0_ports_rsp_payload_data[511:0] ), //i
    .sram_1_ports_cmd_valid         (iCache_1_sram_1_ports_cmd_valid                  ), //o
    .sram_1_ports_cmd_payload_addr  (iCache_1_sram_1_ports_cmd_payload_addr[3:0]      ), //o
    .sram_1_ports_cmd_payload_wen   (iCache_1_sram_1_ports_cmd_payload_wen[15:0]      ), //o
    .sram_1_ports_cmd_payload_wdata (iCache_1_sram_1_ports_cmd_payload_wdata[511:0]   ), //o
    .sram_1_ports_cmd_payload_wstrb (iCache_1_sram_1_ports_cmd_payload_wstrb[63:0]    ), //o
    .sram_1_ports_rsp_valid         (sramBanks_2_sram_1_ports_rsp_valid               ), //i
    .sram_1_ports_rsp_payload_data  (sramBanks_2_sram_1_ports_rsp_payload_data[511:0] ), //i
    .sram_2_ports_cmd_valid         (iCache_1_sram_2_ports_cmd_valid                  ), //o
    .sram_2_ports_cmd_payload_addr  (iCache_1_sram_2_ports_cmd_payload_addr[3:0]      ), //o
    .sram_2_ports_cmd_payload_wen   (iCache_1_sram_2_ports_cmd_payload_wen[15:0]      ), //o
    .sram_2_ports_cmd_payload_wdata (iCache_1_sram_2_ports_cmd_payload_wdata[511:0]   ), //o
    .sram_2_ports_cmd_payload_wstrb (iCache_1_sram_2_ports_cmd_payload_wstrb[63:0]    ), //o
    .sram_2_ports_rsp_valid         (sramBanks_2_sram_2_ports_rsp_valid               ), //i
    .sram_2_ports_rsp_payload_data  (sramBanks_2_sram_2_ports_rsp_payload_data[511:0] ), //i
    .sram_3_ports_cmd_valid         (iCache_1_sram_3_ports_cmd_valid                  ), //o
    .sram_3_ports_cmd_payload_addr  (iCache_1_sram_3_ports_cmd_payload_addr[3:0]      ), //o
    .sram_3_ports_cmd_payload_wen   (iCache_1_sram_3_ports_cmd_payload_wen[15:0]      ), //o
    .sram_3_ports_cmd_payload_wdata (iCache_1_sram_3_ports_cmd_payload_wdata[511:0]   ), //o
    .sram_3_ports_cmd_payload_wstrb (iCache_1_sram_3_ports_cmd_payload_wstrb[63:0]    ), //o
    .sram_3_ports_rsp_valid         (sramBanks_2_sram_3_ports_rsp_valid               ), //i
    .sram_3_ports_rsp_payload_data  (sramBanks_2_sram_3_ports_rsp_payload_data[511:0] ), //i
    .next_level_cmd_valid           (iCache_1_next_level_cmd_valid                    ), //o
    .next_level_cmd_ready           (icache_ar_ready                                  ), //i
    .next_level_cmd_payload_addr    (iCache_1_next_level_cmd_payload_addr[63:0]       ), //o
    .next_level_cmd_payload_len     (iCache_1_next_level_cmd_payload_len[3:0]         ), //o
    .next_level_cmd_payload_size    (iCache_1_next_level_cmd_payload_size[2:0]        ), //o
    .next_level_rsp_valid           (iCache_1_next_level_rsp_valid                    ), //i
    .next_level_rsp_payload_data    (icache_r_payload_data[63:0]                      ), //i
    .io_axiClk                      (io_axiClk                                        ), //i
    .resetCtrl_axiReset             (resetCtrl_axiReset                               )  //i
  );
  SramBanks sramBanks_2 (
    .sram_0_ports_cmd_valid         (iCache_1_sram_0_ports_cmd_valid                 ), //i
    .sram_0_ports_cmd_payload_addr  (iCache_1_sram_0_ports_cmd_payload_addr[3:0]     ), //i
    .sram_0_ports_cmd_payload_wen   (iCache_1_sram_0_ports_cmd_payload_wen[15:0]     ), //i
    .sram_0_ports_cmd_payload_wdata (iCache_1_sram_0_ports_cmd_payload_wdata[511:0]  ), //i
    .sram_0_ports_cmd_payload_wstrb (iCache_1_sram_0_ports_cmd_payload_wstrb[63:0]   ), //i
    .sram_0_ports_rsp_valid         (sramBanks_2_sram_0_ports_rsp_valid              ), //o
    .sram_0_ports_rsp_payload_data  (sramBanks_2_sram_0_ports_rsp_payload_data[511:0]), //o
    .sram_1_ports_cmd_valid         (iCache_1_sram_1_ports_cmd_valid                 ), //i
    .sram_1_ports_cmd_payload_addr  (iCache_1_sram_1_ports_cmd_payload_addr[3:0]     ), //i
    .sram_1_ports_cmd_payload_wen   (iCache_1_sram_1_ports_cmd_payload_wen[15:0]     ), //i
    .sram_1_ports_cmd_payload_wdata (iCache_1_sram_1_ports_cmd_payload_wdata[511:0]  ), //i
    .sram_1_ports_cmd_payload_wstrb (iCache_1_sram_1_ports_cmd_payload_wstrb[63:0]   ), //i
    .sram_1_ports_rsp_valid         (sramBanks_2_sram_1_ports_rsp_valid              ), //o
    .sram_1_ports_rsp_payload_data  (sramBanks_2_sram_1_ports_rsp_payload_data[511:0]), //o
    .sram_2_ports_cmd_valid         (iCache_1_sram_2_ports_cmd_valid                 ), //i
    .sram_2_ports_cmd_payload_addr  (iCache_1_sram_2_ports_cmd_payload_addr[3:0]     ), //i
    .sram_2_ports_cmd_payload_wen   (iCache_1_sram_2_ports_cmd_payload_wen[15:0]     ), //i
    .sram_2_ports_cmd_payload_wdata (iCache_1_sram_2_ports_cmd_payload_wdata[511:0]  ), //i
    .sram_2_ports_cmd_payload_wstrb (iCache_1_sram_2_ports_cmd_payload_wstrb[63:0]   ), //i
    .sram_2_ports_rsp_valid         (sramBanks_2_sram_2_ports_rsp_valid              ), //o
    .sram_2_ports_rsp_payload_data  (sramBanks_2_sram_2_ports_rsp_payload_data[511:0]), //o
    .sram_3_ports_cmd_valid         (iCache_1_sram_3_ports_cmd_valid                 ), //i
    .sram_3_ports_cmd_payload_addr  (iCache_1_sram_3_ports_cmd_payload_addr[3:0]     ), //i
    .sram_3_ports_cmd_payload_wen   (iCache_1_sram_3_ports_cmd_payload_wen[15:0]     ), //i
    .sram_3_ports_cmd_payload_wdata (iCache_1_sram_3_ports_cmd_payload_wdata[511:0]  ), //i
    .sram_3_ports_cmd_payload_wstrb (iCache_1_sram_3_ports_cmd_payload_wstrb[63:0]   ), //i
    .sram_3_ports_rsp_valid         (sramBanks_2_sram_3_ports_rsp_valid              ), //o
    .sram_3_ports_rsp_payload_data  (sramBanks_2_sram_3_ports_rsp_payload_data[511:0]), //o
    .io_axiClk                      (io_axiClk                                       ), //i
    .resetCtrl_axiReset             (resetCtrl_axiReset                              )  //i
  );
  DCache dCache_1 (
    .stall                          (dCache_1_stall                                    ), //o
    .flush                          (1'b0                                              ), //i
    .cpu_cmd_valid                  (DCachePlugin_dcache_access_cmd_valid              ), //i
    .cpu_cmd_ready                  (dCache_1_cpu_cmd_ready                            ), //o
    .cpu_cmd_payload_addr           (DCachePlugin_dcache_access_cmd_payload_addr[63:0] ), //i
    .cpu_cmd_payload_wen            (DCachePlugin_dcache_access_cmd_payload_wen        ), //i
    .cpu_cmd_payload_wdata          (DCachePlugin_dcache_access_cmd_payload_wdata[63:0]), //i
    .cpu_cmd_payload_wstrb          (DCachePlugin_dcache_access_cmd_payload_wstrb[7:0] ), //i
    .cpu_cmd_payload_size           (DCachePlugin_dcache_access_cmd_payload_size[2:0]  ), //i
    .cpu_rsp_valid                  (dCache_1_cpu_rsp_valid                            ), //o
    .cpu_rsp_payload_data           (dCache_1_cpu_rsp_payload_data[63:0]               ), //o
    .sram_0_ports_cmd_valid         (dCache_1_sram_0_ports_cmd_valid                   ), //o
    .sram_0_ports_cmd_payload_addr  (dCache_1_sram_0_ports_cmd_payload_addr[1:0]       ), //o
    .sram_0_ports_cmd_payload_wen   (dCache_1_sram_0_ports_cmd_payload_wen[7:0]        ), //o
    .sram_0_ports_cmd_payload_wdata (dCache_1_sram_0_ports_cmd_payload_wdata[511:0]    ), //o
    .sram_0_ports_cmd_payload_wstrb (dCache_1_sram_0_ports_cmd_payload_wstrb[63:0]     ), //o
    .sram_0_ports_rsp_valid         (sramBanks_3_sram_0_ports_rsp_valid                ), //i
    .sram_0_ports_rsp_payload_data  (sramBanks_3_sram_0_ports_rsp_payload_data[511:0]  ), //i
    .sram_1_ports_cmd_valid         (dCache_1_sram_1_ports_cmd_valid                   ), //o
    .sram_1_ports_cmd_payload_addr  (dCache_1_sram_1_ports_cmd_payload_addr[1:0]       ), //o
    .sram_1_ports_cmd_payload_wen   (dCache_1_sram_1_ports_cmd_payload_wen[7:0]        ), //o
    .sram_1_ports_cmd_payload_wdata (dCache_1_sram_1_ports_cmd_payload_wdata[511:0]    ), //o
    .sram_1_ports_cmd_payload_wstrb (dCache_1_sram_1_ports_cmd_payload_wstrb[63:0]     ), //o
    .sram_1_ports_rsp_valid         (sramBanks_3_sram_1_ports_rsp_valid                ), //i
    .sram_1_ports_rsp_payload_data  (sramBanks_3_sram_1_ports_rsp_payload_data[511:0]  ), //i
    .sram_2_ports_cmd_valid         (dCache_1_sram_2_ports_cmd_valid                   ), //o
    .sram_2_ports_cmd_payload_addr  (dCache_1_sram_2_ports_cmd_payload_addr[1:0]       ), //o
    .sram_2_ports_cmd_payload_wen   (dCache_1_sram_2_ports_cmd_payload_wen[7:0]        ), //o
    .sram_2_ports_cmd_payload_wdata (dCache_1_sram_2_ports_cmd_payload_wdata[511:0]    ), //o
    .sram_2_ports_cmd_payload_wstrb (dCache_1_sram_2_ports_cmd_payload_wstrb[63:0]     ), //o
    .sram_2_ports_rsp_valid         (sramBanks_3_sram_2_ports_rsp_valid                ), //i
    .sram_2_ports_rsp_payload_data  (sramBanks_3_sram_2_ports_rsp_payload_data[511:0]  ), //i
    .sram_3_ports_cmd_valid         (dCache_1_sram_3_ports_cmd_valid                   ), //o
    .sram_3_ports_cmd_payload_addr  (dCache_1_sram_3_ports_cmd_payload_addr[1:0]       ), //o
    .sram_3_ports_cmd_payload_wen   (dCache_1_sram_3_ports_cmd_payload_wen[7:0]        ), //o
    .sram_3_ports_cmd_payload_wdata (dCache_1_sram_3_ports_cmd_payload_wdata[511:0]    ), //o
    .sram_3_ports_cmd_payload_wstrb (dCache_1_sram_3_ports_cmd_payload_wstrb[63:0]     ), //o
    .sram_3_ports_rsp_valid         (sramBanks_3_sram_3_ports_rsp_valid                ), //i
    .sram_3_ports_rsp_payload_data  (sramBanks_3_sram_3_ports_rsp_payload_data[511:0]  ), //i
    .next_level_cmd_valid           (dCache_1_next_level_cmd_valid                     ), //o
    .next_level_cmd_ready           (1'b1                                              ), //i
    .next_level_cmd_payload_addr    (dCache_1_next_level_cmd_payload_addr[63:0]        ), //o
    .next_level_cmd_payload_len     (dCache_1_next_level_cmd_payload_len[3:0]          ), //o
    .next_level_cmd_payload_size    (dCache_1_next_level_cmd_payload_size[2:0]         ), //o
    .next_level_cmd_payload_wen     (dCache_1_next_level_cmd_payload_wen               ), //o
    .next_level_cmd_payload_wdata   (dCache_1_next_level_cmd_payload_wdata[63:0]       ), //o
    .next_level_cmd_payload_wstrb   (dCache_1_next_level_cmd_payload_wstrb[7:0]        ), //o
    .next_level_rsp_valid           (dCache_1_next_level_rsp_valid                     ), //i
    .next_level_rsp_payload_data    (dcache_r_payload_data[63:0]                       ), //i
    .next_level_rsp_payload_bresp   (dcache_b_payload_resp[1:0]                        ), //i
    .next_level_rsp_payload_rvalid  (dCache_1_next_level_rsp_payload_rvalid            ), //i
    .cpu_bypass_cmd_valid           (dCache_1_cpu_bypass_cmd_valid                     ), //o
    .cpu_bypass_cmd_ready           (1'b1                                              ), //i
    .cpu_bypass_cmd_payload_addr    (dCache_1_cpu_bypass_cmd_payload_addr[63:0]        ), //o
    .cpu_bypass_cmd_payload_wen     (dCache_1_cpu_bypass_cmd_payload_wen               ), //o
    .cpu_bypass_cmd_payload_wdata   (dCache_1_cpu_bypass_cmd_payload_wdata[63:0]       ), //o
    .cpu_bypass_cmd_payload_wstrb   (dCache_1_cpu_bypass_cmd_payload_wstrb[7:0]        ), //o
    .cpu_bypass_cmd_payload_size    (dCache_1_cpu_bypass_cmd_payload_size[2:0]         ), //o
    .cpu_bypass_rsp_valid           (dCache_1_cpu_bypass_rsp_valid                     ), //i
    .cpu_bypass_rsp_payload_data    (dcache_r_payload_data[63:0]                       ), //i
    .io_axiClk                      (io_axiClk                                         ), //i
    .resetCtrl_axiReset             (resetCtrl_axiReset                                )  //i
  );
  SramBanks_1 sramBanks_3 (
    .sram_0_ports_cmd_valid         (dCache_1_sram_0_ports_cmd_valid                 ), //i
    .sram_0_ports_cmd_payload_addr  (dCache_1_sram_0_ports_cmd_payload_addr[1:0]     ), //i
    .sram_0_ports_cmd_payload_wen   (dCache_1_sram_0_ports_cmd_payload_wen[7:0]      ), //i
    .sram_0_ports_cmd_payload_wdata (dCache_1_sram_0_ports_cmd_payload_wdata[511:0]  ), //i
    .sram_0_ports_cmd_payload_wstrb (dCache_1_sram_0_ports_cmd_payload_wstrb[63:0]   ), //i
    .sram_0_ports_rsp_valid         (sramBanks_3_sram_0_ports_rsp_valid              ), //o
    .sram_0_ports_rsp_payload_data  (sramBanks_3_sram_0_ports_rsp_payload_data[511:0]), //o
    .sram_1_ports_cmd_valid         (dCache_1_sram_1_ports_cmd_valid                 ), //i
    .sram_1_ports_cmd_payload_addr  (dCache_1_sram_1_ports_cmd_payload_addr[1:0]     ), //i
    .sram_1_ports_cmd_payload_wen   (dCache_1_sram_1_ports_cmd_payload_wen[7:0]      ), //i
    .sram_1_ports_cmd_payload_wdata (dCache_1_sram_1_ports_cmd_payload_wdata[511:0]  ), //i
    .sram_1_ports_cmd_payload_wstrb (dCache_1_sram_1_ports_cmd_payload_wstrb[63:0]   ), //i
    .sram_1_ports_rsp_valid         (sramBanks_3_sram_1_ports_rsp_valid              ), //o
    .sram_1_ports_rsp_payload_data  (sramBanks_3_sram_1_ports_rsp_payload_data[511:0]), //o
    .sram_2_ports_cmd_valid         (dCache_1_sram_2_ports_cmd_valid                 ), //i
    .sram_2_ports_cmd_payload_addr  (dCache_1_sram_2_ports_cmd_payload_addr[1:0]     ), //i
    .sram_2_ports_cmd_payload_wen   (dCache_1_sram_2_ports_cmd_payload_wen[7:0]      ), //i
    .sram_2_ports_cmd_payload_wdata (dCache_1_sram_2_ports_cmd_payload_wdata[511:0]  ), //i
    .sram_2_ports_cmd_payload_wstrb (dCache_1_sram_2_ports_cmd_payload_wstrb[63:0]   ), //i
    .sram_2_ports_rsp_valid         (sramBanks_3_sram_2_ports_rsp_valid              ), //o
    .sram_2_ports_rsp_payload_data  (sramBanks_3_sram_2_ports_rsp_payload_data[511:0]), //o
    .sram_3_ports_cmd_valid         (dCache_1_sram_3_ports_cmd_valid                 ), //i
    .sram_3_ports_cmd_payload_addr  (dCache_1_sram_3_ports_cmd_payload_addr[1:0]     ), //i
    .sram_3_ports_cmd_payload_wen   (dCache_1_sram_3_ports_cmd_payload_wen[7:0]      ), //i
    .sram_3_ports_cmd_payload_wdata (dCache_1_sram_3_ports_cmd_payload_wdata[511:0]  ), //i
    .sram_3_ports_cmd_payload_wstrb (dCache_1_sram_3_ports_cmd_payload_wstrb[63:0]   ), //i
    .sram_3_ports_rsp_valid         (sramBanks_3_sram_3_ports_rsp_valid              ), //o
    .sram_3_ports_rsp_payload_data  (sramBanks_3_sram_3_ports_rsp_payload_data[511:0]), //o
    .io_axiClk                      (io_axiClk                                       ), //i
    .resetCtrl_axiReset             (resetCtrl_axiReset                              )  //i
  );
  assign writeback_RD = (writeback_IS_LOAD ? writeback_LSU_RDATA : writeback_ALU_RESULT);
  assign memaccess_LSU_HOLD = DCachePlugin_dcache_access_stall;
  assign memaccess_TIMER_CEN = ((memaccess_LSUPlugin_is_timer && memaccess_LSUPlugin_is_mem) && memaccess_arbitration_isFiring);
  assign memaccess_LSU_WDATA = memaccess_LSUPlugin_lsu_wdata;
  assign execute_INT_HOLD = clint_1_int_hold;
  assign execute_REDIRECT_PC_NEXT = execute_ALUPlugin_redirect_pc_next;
  assign execute_REDIRECT_VALID = execute_ALUPlugin_redirect_valid;
  assign execute_IS_RET = execute_ALUPlugin_is_ret;
  assign execute_IS_CALL = execute_ALUPlugin_is_call;
  assign execute_IS_JMP = execute_ALUPlugin_is_jmp;
  assign execute_BRANCH_HISTORY = execute_ALUPlugin_branch_history;
  assign execute_BRANCH_TAKEN = execute_ALUPlugin_branch_taken;
  assign execute_BRANCH_OR_JUMP = (execute_ALUPlugin_branch_or_jump && execute_arbitration_isFiring);
  assign execute_BRANCH_OR_JALR = execute_ALUPlugin_branch_or_jalr;
  assign execute_MEM_WDATA = (execute_RS2_FROM_WB ? _zz_execute_MEM_WDATA_2 : (execute_RS2_FROM_MEM ? _zz_execute_MEM_WDATA_1 : (execute_RS2_FROM_LOAD ? _zz_execute_MEM_WDATA : execute_RS2)));
  assign execute_ALU_RESULT = execute_ALUPlugin_alu_result;
  assign decode_CSR_RDATA = csrRegfile_1_cpu_ports_rdata;
  assign execute_CSR_WEN = decode_to_execute_CSR_WEN;
  assign decode_CSR_WEN = decode_DecodePlugin_csr_wen;
  assign execute_CSR_ADDR = decode_to_execute_CSR_ADDR;
  assign decode_CSR_ADDR = decode_DecodePlugin_csr_addr;
  assign decode_CSR_CTRL = decode_DecodePlugin_csr_ctrl;
  assign execute_IS_STORE = decode_to_execute_IS_STORE;
  assign decode_IS_STORE = decode_DecodePlugin_is_store;
  assign execute_IS_LOAD = decode_to_execute_IS_LOAD;
  assign decode_IS_LOAD = decode_DecodePlugin_is_load;
  assign writeback_RD_ADDR = memaccess_to_writeback_RD_ADDR;
  assign memaccess_RD_ADDR = execute_to_memaccess_RD_ADDR;
  assign decode_RD_ADDR = decode_DecodePlugin_rd_addr;
  assign writeback_RD_WEN = memaccess_to_writeback_RD_WEN;
  assign memaccess_RD_WEN = execute_to_memaccess_RD_WEN;
  assign execute_RD_WEN = decode_to_execute_RD_WEN;
  assign decode_RD_WEN = decode_DecodePlugin_rd_wen;
  assign execute_MEM_CTRL = decode_to_execute_MEM_CTRL;
  assign decode_MEM_CTRL = decode_DecodePlugin_mem_ctrl;
  assign decode_SRC2_IS_IMM = decode_DecodePlugin_src2_is_imm;
  assign decode_ALU_WORD = decode_DecodePlugin_alu_word;
  assign decode_ALU_CTRL = decode_DecodePlugin_alu_ctrl;
  assign execute_RS2_ADDR = decode_to_execute_RS2_ADDR;
  assign decode_RS2_ADDR = decode_DecodePlugin_rs2_addr;
  assign decode_RS1_ADDR = decode_DecodePlugin_rs1_addr;
  assign decode_RS2 = decode_DecodePlugin_rs2;
  assign decode_RS1 = decode_DecodePlugin_rs1;
  assign decode_IMM = decode_DecodePlugin_imm;
  assign fetch_INT_PC = clint_1_int_pc;
  assign fetch_INT_EN = clint_1_int_en;
  assign fetch_PREDICT_PC = pc_next;
  assign decode_PREDICT_TAKEN = fetch_to_decode_PREDICT_TAKEN;
  assign fetch_PREDICT_TAKEN = fetch_FetchPlugin_predict_taken_out_payload;
  assign fetch_PREDICT_VALID = ICachePlugin_icache_access_cmd_fire_4;
  assign memaccess_INSTRUCTION = execute_to_memaccess_INSTRUCTION;
  assign execute_INSTRUCTION = decode_to_execute_INSTRUCTION;
  assign fetch_INSTRUCTION = fetch_FetchPlugin_instruction_out_stream_payload;
  assign decode_PC_NEXT = fetch_to_decode_PC_NEXT;
  assign fetch_PC_NEXT = fetch_FetchPlugin_pc_stream_fifo_next_payload;
  assign memaccess_PC = execute_to_memaccess_PC;
  assign fetch_PC = fetch_FetchPlugin_pc_out_stream_payload;
  assign writeback_INSTRUCTION = memaccess_to_writeback_INSTRUCTION;
  assign writeback_PC = memaccess_to_writeback_PC;
  assign writeback_ALU_RESULT = memaccess_to_writeback_ALU_RESULT;
  assign writeback_LSU_RDATA = memaccess_to_writeback_LSU_RDATA;
  assign writeback_IS_LOAD = memaccess_to_writeback_IS_LOAD;
  assign memaccess_MEM_CTRL = execute_to_memaccess_MEM_CTRL;
  assign memaccess_MEM_WDATA = execute_to_memaccess_MEM_WDATA;
  assign memaccess_IS_STORE = execute_to_memaccess_IS_STORE;
  assign memaccess_IS_LOAD = execute_to_memaccess_IS_LOAD;
  assign execute_CSR_CTRL = decode_to_execute_CSR_CTRL;
  assign execute_SRC1 = execute_ALUPlugin_src1;
  assign _zz_ecall = execute_CSR_CTRL;
  assign _zz_decode_to_execute_CSR_ADDR = decode_CSR_ADDR;
  assign _zz_memaccess_arbitration_haltItself = memaccess_LSU_HOLD;
  assign _zz_DecodePlugin_hazard_ctrl_rs1_from_mem = execute_BRANCH_OR_JALR;
  assign _zz_DecodePlugin_hazard_rs2_from_mem = execute_RS2_ADDR;
  assign _zz_DecodePlugin_hazard_rs1_from_mem = memaccess_IS_LOAD;
  assign _zz_DecodePlugin_hazard_rs1_from_mem_1 = execute_RS1_ADDR;
  assign _zz_DecodePlugin_hazard_rs1_from_mem_2 = memaccess_RD_ADDR;
  assign _zz_DecodePlugin_hazard_rs1_from_mem_3 = memaccess_RD_WEN;
  assign execute_PC_NEXT = decode_to_execute_PC_NEXT;
  assign execute_PREDICT_TAKEN = decode_to_execute_PREDICT_TAKEN;
  assign execute_CSR_RDATA = decode_to_execute_CSR_RDATA;
  assign execute_ALU_WORD = decode_to_execute_ALU_WORD;
  assign execute_CTRL_RS2_FROM_WB = DecodePlugin_hazard_ctrl_rs2_from_wb;
  assign execute_CTRL_RS2_FROM_LOAD = DecodePlugin_hazard_ctrl_rs2_from_load;
  assign execute_CTRL_RS2_FROM_MEM = DecodePlugin_hazard_ctrl_rs2_from_mem;
  assign execute_CTRL_RS1_FROM_WB = DecodePlugin_hazard_ctrl_rs1_from_wb;
  assign _zz_execute_MEM_WDATA = memaccess_LSU_RDATA;
  assign execute_CTRL_RS1_FROM_LOAD = DecodePlugin_hazard_ctrl_rs1_from_load;
  assign _zz_execute_MEM_WDATA_1 = memaccess_ALU_RESULT;
  assign execute_CTRL_RS1_FROM_MEM = DecodePlugin_hazard_ctrl_rs1_from_mem;
  assign execute_RS2 = decode_to_execute_RS2;
  assign execute_RS2_FROM_WB = DecodePlugin_hazard_rs2_from_wb;
  assign execute_RS2_FROM_LOAD = DecodePlugin_hazard_rs2_from_load;
  assign execute_RS2_FROM_MEM = DecodePlugin_hazard_rs2_from_mem;
  assign execute_IMM = decode_to_execute_IMM;
  assign execute_SRC2_IS_IMM = decode_to_execute_SRC2_IS_IMM;
  assign execute_RS1 = decode_to_execute_RS1;
  assign execute_RS1_FROM_WB = DecodePlugin_hazard_rs1_from_wb;
  assign memaccess_LSU_RDATA = memaccess_LSUPlugin_lsu_rdata;
  assign execute_RS1_FROM_LOAD = DecodePlugin_hazard_rs1_from_load;
  assign memaccess_ALU_RESULT = execute_to_memaccess_ALU_RESULT;
  assign execute_RS1_FROM_MEM = DecodePlugin_hazard_rs1_from_mem;
  assign execute_PC = decode_to_execute_PC;
  assign execute_RS1_ADDR = decode_to_execute_RS1_ADDR;
  assign execute_RD_ADDR = decode_to_execute_RD_ADDR;
  assign execute_ALU_CTRL = decode_to_execute_ALU_CTRL;
  assign _zz_execute_MEM_WDATA_2 = writeback_RD;
  assign _zz_DecodePlugin_hazard_rs1_from_wb = writeback_RD_ADDR;
  assign _zz_DecodePlugin_hazard_rs1_from_wb_1 = writeback_RD_WEN;
  assign decode_INSTRUCTION = fetch_to_decode_INSTRUCTION;
  assign decode_PC = fetch_to_decode_PC;
  assign _zz_execute_to_memaccess_PC = execute_PC;
  assign fetch_BPU_PC_NEXT = gshare_predictor_1_predict_pc_next;
  assign _zz_pc_next = execute_REDIRECT_PC_NEXT;
  assign when_FetchPlugin_l97 = execute_REDIRECT_VALID;
  assign fetch_BPU_BRANCH_TAKEN = gshare_predictor_1_predict_taken;
  assign when_FetchPlugin_l94 = fetch_INT_EN;
  assign fetch_arbitration_haltByOther = 1'b0;
  always @(*) begin
    fetch_arbitration_removeIt = 1'b0;
    if(fetch_arbitration_isFlushed) begin
      fetch_arbitration_removeIt = 1'b1;
    end
  end

  assign fetch_arbitration_flushNext = 1'b0;
  assign decode_arbitration_haltByOther = 1'b0;
  always @(*) begin
    decode_arbitration_removeIt = 1'b0;
    if(decode_arbitration_isFlushed) begin
      decode_arbitration_removeIt = 1'b1;
    end
  end

  assign decode_arbitration_flushNext = 1'b0;
  assign execute_arbitration_haltByOther = 1'b0;
  always @(*) begin
    execute_arbitration_removeIt = 1'b0;
    if(execute_arbitration_isFlushed) begin
      execute_arbitration_removeIt = 1'b1;
    end
  end

  assign execute_arbitration_flushNext = 1'b0;
  assign memaccess_arbitration_haltByOther = 1'b0;
  always @(*) begin
    memaccess_arbitration_removeIt = 1'b0;
    if(memaccess_arbitration_isFlushed) begin
      memaccess_arbitration_removeIt = 1'b1;
    end
  end

  assign memaccess_arbitration_flushNext = 1'b0;
  assign writeback_arbitration_haltByOther = 1'b0;
  always @(*) begin
    writeback_arbitration_removeIt = 1'b0;
    if(writeback_arbitration_isFlushed) begin
      writeback_arbitration_removeIt = 1'b1;
    end
  end

  assign writeback_arbitration_flushNext = 1'b0;
  assign fetch_FetchPlugin_fetch_flush = (when_FetchPlugin_l94 || fetch_arbitration_flushIt);
  assign ICachePlugin_icache_access_cmd_fire = (ICachePlugin_icache_access_cmd_valid && ICachePlugin_icache_access_cmd_ready);
  assign fetch_FetchPlugin_bpu_predict_taken = (fetch_BPU_BRANCH_TAKEN && ICachePlugin_icache_access_cmd_fire);
  assign fetch_FetchPlugin_fifo_all_valid = ((fetch_FetchPlugin_pc_out_stream_valid && fetch_FetchPlugin_instruction_out_stream_valid) && fetch_FetchPlugin_pc_stream_fifo_next_valid);
  assign IDLE = 2'b00;
  assign FETCH = 2'b01;
  assign HALT = 2'b11;
  assign when_FetchPlugin_l64 = (! fetch_arbitration_isStuck);
  always @(*) begin
    if((fetch_state == IDLE)) begin
        if(when_FetchPlugin_l64) begin
          fetch_state_next = FETCH;
        end else begin
          fetch_state_next = IDLE;
        end
    end else if((fetch_state == FETCH)) begin
        if(when_FetchPlugin_l72) begin
          fetch_state_next = HALT;
        end else begin
          fetch_state_next = FETCH;
        end
    end else if((fetch_state == HALT)) begin
        if(when_FetchPlugin_l80) begin
          fetch_state_next = FETCH;
        end else begin
          fetch_state_next = HALT;
        end
    end else begin
        fetch_state_next = IDLE;
    end
  end

  assign ICachePlugin_icache_access_cmd_isStall = (ICachePlugin_icache_access_cmd_valid && (! ICachePlugin_icache_access_cmd_ready));
  assign when_FetchPlugin_l72 = (ICachePlugin_icache_access_cmd_isStall || fetch_arbitration_isStuck);
  assign when_FetchPlugin_l80 = (ICachePlugin_icache_access_cmd_ready && (! fetch_arbitration_isStuck));
  assign when_FetchPlugin_l93 = (! ICachePlugin_icache_access_cmd_ready);
  assign when_FetchPlugin_l109 = (fetch_state_next == FETCH);
  assign ICachePlugin_icache_access_cmd_fire_1 = (ICachePlugin_icache_access_cmd_valid && ICachePlugin_icache_access_cmd_ready);
  assign ICachePlugin_icache_access_cmd_fire_2 = (ICachePlugin_icache_access_cmd_valid && ICachePlugin_icache_access_cmd_ready);
  assign fetch_FetchPlugin_pc_in_stream_valid = ICachePlugin_icache_access_cmd_fire_2;
  assign fetch_FetchPlugin_pc_in_stream_payload = pc_next;
  assign fetch_FetchPlugin_pc_out_stream_ready = fetch_arbitration_isFiring;
  assign fetch_FetchPlugin_pc_in_stream_ready = fetch_FetchPlugin_pc_stream_fifo_ports_s_ports_ready;
  assign fetch_FetchPlugin_pc_out_stream_valid = fetch_FetchPlugin_pc_stream_fifo_ports_m_ports_valid;
  assign fetch_FetchPlugin_pc_out_stream_payload = fetch_FetchPlugin_pc_stream_fifo_ports_m_ports_payload;
  assign ICachePlugin_icache_access_cmd_fire_3 = (ICachePlugin_icache_access_cmd_valid && ICachePlugin_icache_access_cmd_ready);
  assign fetch_FetchPlugin_predict_taken_in_valid = ICachePlugin_icache_access_cmd_fire_3;
  assign fetch_FetchPlugin_predict_taken_in_payload = fetch_BPU_BRANCH_TAKEN;
  assign fetch_FetchPlugin_predict_taken_out_ready = fetch_arbitration_isFiring;
  assign fetch_FetchPlugin_predict_taken_in_ready = fetch_FetchPlugin_predict_taken_fifo_ports_s_ports_ready;
  assign fetch_FetchPlugin_predict_taken_out_valid = fetch_FetchPlugin_predict_taken_fifo_ports_m_ports_valid;
  assign fetch_FetchPlugin_predict_taken_out_payload = fetch_FetchPlugin_predict_taken_fifo_ports_m_ports_payload;
  assign fetch_FetchPlugin_instruction_in_stream_valid = ((ICachePlugin_icache_access_rsp_valid && (! rsp_flush)) && (! fetch_FetchPlugin_fetch_flush));
  assign fetch_FetchPlugin_instruction_in_stream_payload = ICachePlugin_icache_access_rsp_payload_data;
  assign fetch_FetchPlugin_instruction_out_stream_ready = fetch_arbitration_isFiring;
  assign fetch_FetchPlugin_instruction_in_stream_ready = fetch_FetchPlugin_instruction_stream_fifo_ports_s_ports_ready;
  assign fetch_FetchPlugin_instruction_out_stream_valid = fetch_FetchPlugin_instruction_stream_fifo_ports_m_ports_valid;
  assign fetch_FetchPlugin_instruction_out_stream_payload = fetch_FetchPlugin_instruction_stream_fifo_ports_m_ports_payload;
  assign ICachePlugin_icache_access_cmd_fire_4 = (ICachePlugin_icache_access_cmd_valid && ICachePlugin_icache_access_cmd_ready);
  assign fetch_arbitration_isValid = ((fetch_FetchPlugin_fifo_all_valid && (! fetch_arbitration_isStuck)) && (! fetch_FetchPlugin_fetch_flush));
  assign ICachePlugin_icache_access_cmd_valid = (fetch_valid && (! fetch_FetchPlugin_fetch_flush));
  assign ICachePlugin_icache_access_cmd_payload_addr = pc_next;
  assign decode_DecodePlugin_rs1_req = (! (((decode_INSTRUCTION[6 : 0] == 7'h37) || (decode_INSTRUCTION[6 : 0] == 7'h17)) || (decode_INSTRUCTION[6 : 0] == 7'h6f)));
  assign decode_DecodePlugin_rs2_req = (! ((((decode_INSTRUCTION[6 : 0] == 7'h37) || (decode_INSTRUCTION[6 : 0] == 7'h17)) || (decode_INSTRUCTION[6 : 0] == 7'h6f)) || ((((decode_INSTRUCTION[6 : 0] == 7'h13) || (decode_INSTRUCTION[6 : 0] == 7'h1b)) || (decode_INSTRUCTION[6 : 0] == 7'h03)) || (decode_INSTRUCTION[6 : 0] == 7'h67))));
  assign decode_DecodePlugin_rs1_addr = decode_INSTRUCTION[19 : 15];
  assign decode_DecodePlugin_rs2_addr = decode_INSTRUCTION[24 : 20];
  assign decode_DecodePlugin_rd_addr = decode_INSTRUCTION[11 : 7];
  assign decode_DecodePlugin_alu_word = ((decode_INSTRUCTION[6 : 0] == 7'h3b) || (decode_INSTRUCTION[6 : 0] == 7'h1b));
  assign decode_DecodePlugin_src2_is_imm = ((((((decode_INSTRUCTION[6 : 0] == 7'h13) || (decode_INSTRUCTION[6 : 0] == 7'h1b)) || (decode_INSTRUCTION[6 : 0] == 7'h03)) || (decode_INSTRUCTION[6 : 0] == 7'h67)) || (decode_INSTRUCTION[6 : 0] == 7'h23)) || ((decode_INSTRUCTION[6 : 0] == 7'h37) || (decode_INSTRUCTION[6 : 0] == 7'h17)));
  assign decode_DecodePlugin_csr_addr = decode_INSTRUCTION[31 : 20];
  assign decode_DecodePlugin_csr_wen = (((decode_DecodePlugin_csr_ctrl == CsrCtrlEnum_CSRRW) || (decode_DecodePlugin_csr_ctrl == CsrCtrlEnum_CSRRS)) || (decode_DecodePlugin_csr_ctrl == CsrCtrlEnum_CSRRC));
  assign when_DecodePlugin_l116 = ((((decode_INSTRUCTION[6 : 0] == 7'h13) || (decode_INSTRUCTION[6 : 0] == 7'h1b)) || (decode_INSTRUCTION[6 : 0] == 7'h03)) || (decode_INSTRUCTION[6 : 0] == 7'h67));
  assign _zz_decode_DecodePlugin_imm = decode_INSTRUCTION[31];
  always @(*) begin
    _zz_decode_DecodePlugin_imm_1[51] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[50] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[49] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[48] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[47] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[46] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[45] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[44] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[43] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[42] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[41] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[40] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[39] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[38] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[37] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[36] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[35] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[34] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[33] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[32] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[31] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[30] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[29] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[28] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[27] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[26] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[25] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[24] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[23] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[22] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[21] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[20] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[19] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[18] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[17] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[16] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[15] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[14] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[13] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[12] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[11] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[10] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[9] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[8] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[7] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[6] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[5] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[4] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[3] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[2] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[1] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[0] = _zz_decode_DecodePlugin_imm;
  end

  always @(*) begin
    if(when_DecodePlugin_l116) begin
      decode_DecodePlugin_imm = {_zz_decode_DecodePlugin_imm_1,decode_INSTRUCTION[31 : 20]};
    end else begin
      if(when_DecodePlugin_l119) begin
        decode_DecodePlugin_imm = {_zz_decode_DecodePlugin_imm_3,{decode_INSTRUCTION[31 : 25],decode_INSTRUCTION[11 : 7]}};
      end else begin
        if(when_DecodePlugin_l122) begin
          decode_DecodePlugin_imm = {{_zz_decode_DecodePlugin_imm_5,{{{decode_INSTRUCTION[31],decode_INSTRUCTION[7]},decode_INSTRUCTION[30 : 25]},decode_INSTRUCTION[11 : 8]}},1'b0};
        end else begin
          if(when_DecodePlugin_l125) begin
            decode_DecodePlugin_imm = {{_zz_decode_DecodePlugin_imm_7,{{{decode_INSTRUCTION[31],decode_INSTRUCTION[19 : 12]},decode_INSTRUCTION[20]},decode_INSTRUCTION[30 : 21]}},1'b0};
          end else begin
            if(when_DecodePlugin_l128) begin
              decode_DecodePlugin_imm = {_zz_decode_DecodePlugin_imm_9,{decode_INSTRUCTION[31 : 12],12'h0}};
            end else begin
              decode_DecodePlugin_imm = {_zz_decode_DecodePlugin_imm_11,decode_INSTRUCTION[31 : 20]};
            end
          end
        end
      end
    end
  end

  assign _zz_decode_DecodePlugin_imm_2 = _zz__zz_decode_DecodePlugin_imm_2[11];
  always @(*) begin
    _zz_decode_DecodePlugin_imm_3[51] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[50] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[49] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[48] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[47] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[46] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[45] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[44] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[43] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[42] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[41] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[40] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[39] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[38] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[37] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[36] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[35] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[34] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[33] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[32] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[31] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[30] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[29] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[28] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[27] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[26] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[25] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[24] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[23] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[22] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[21] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[20] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[19] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[18] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[17] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[16] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[15] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[14] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[13] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[12] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[11] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[10] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[9] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[8] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[7] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[6] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[5] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[4] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[3] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[2] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[1] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[0] = _zz_decode_DecodePlugin_imm_2;
  end

  assign _zz_decode_DecodePlugin_imm_4 = _zz__zz_decode_DecodePlugin_imm_4[11];
  always @(*) begin
    _zz_decode_DecodePlugin_imm_5[50] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[49] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[48] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[47] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[46] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[45] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[44] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[43] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[42] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[41] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[40] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[39] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[38] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[37] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[36] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[35] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[34] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[33] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[32] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[31] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[30] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[29] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[28] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[27] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[26] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[25] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[24] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[23] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[22] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[21] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[20] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[19] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[18] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[17] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[16] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[15] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[14] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[13] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[12] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[11] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[10] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[9] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[8] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[7] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[6] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[5] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[4] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[3] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[2] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[1] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[0] = _zz_decode_DecodePlugin_imm_4;
  end

  assign _zz_decode_DecodePlugin_imm_6 = _zz__zz_decode_DecodePlugin_imm_6[19];
  always @(*) begin
    _zz_decode_DecodePlugin_imm_7[42] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[41] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[40] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[39] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[38] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[37] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[36] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[35] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[34] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[33] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[32] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[31] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[30] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[29] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[28] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[27] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[26] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[25] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[24] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[23] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[22] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[21] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[20] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[19] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[18] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[17] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[16] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[15] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[14] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[13] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[12] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[11] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[10] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[9] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[8] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[7] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[6] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[5] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[4] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[3] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[2] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[1] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[0] = _zz_decode_DecodePlugin_imm_6;
  end

  assign _zz_decode_DecodePlugin_imm_8 = _zz__zz_decode_DecodePlugin_imm_8[31];
  always @(*) begin
    _zz_decode_DecodePlugin_imm_9[31] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[30] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[29] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[28] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[27] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[26] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[25] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[24] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[23] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[22] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[21] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[20] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[19] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[18] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[17] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[16] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[15] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[14] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[13] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[12] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[11] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[10] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[9] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[8] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[7] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[6] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[5] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[4] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[3] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[2] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[1] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[0] = _zz_decode_DecodePlugin_imm_8;
  end

  assign _zz_decode_DecodePlugin_imm_10 = decode_INSTRUCTION[31];
  always @(*) begin
    _zz_decode_DecodePlugin_imm_11[51] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[50] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[49] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[48] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[47] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[46] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[45] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[44] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[43] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[42] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[41] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[40] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[39] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[38] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[37] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[36] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[35] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[34] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[33] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[32] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[31] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[30] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[29] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[28] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[27] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[26] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[25] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[24] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[23] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[22] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[21] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[20] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[19] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[18] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[17] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[16] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[15] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[14] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[13] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[12] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[11] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[10] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[9] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[8] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[7] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[6] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[5] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[4] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[3] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[2] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[1] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[0] = _zz_decode_DecodePlugin_imm_10;
  end

  assign when_DecodePlugin_l119 = (decode_INSTRUCTION[6 : 0] == 7'h23);
  assign when_DecodePlugin_l122 = (decode_INSTRUCTION[6 : 0] == 7'h63);
  assign when_DecodePlugin_l125 = (decode_INSTRUCTION[6 : 0] == 7'h6f);
  assign when_DecodePlugin_l128 = ((decode_INSTRUCTION[6 : 0] == 7'h37) || (decode_INSTRUCTION[6 : 0] == 7'h17));
  always @(*) begin
    casez(decode_INSTRUCTION)
      32'b0000000??????????000?????0110011, 32'b0000000??????????000?????0111011, 32'b?????????????????000?????0010011, 32'b?????????????????000?????0011011, 32'b?????????????????000?????0100011, 32'b?????????????????001?????0100011, 32'b?????????????????010?????0100011, 32'b?????????????????011?????0100011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_ADD;
      end
      32'b0100000??????????000?????0110011, 32'b0100000??????????000?????0111011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_SUB;
      end
      32'b0000000??????????010?????0110011, 32'b?????????????????010?????0010011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_SLT;
      end
      32'b0000000??????????011?????0110011, 32'b?????????????????011?????0010011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_SLTU;
      end
      32'b0000000??????????100?????0110011, 32'b?????????????????100?????0010011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_XOR_1;
      end
      32'b0000000??????????001?????0110011, 32'b000000???????????001?????0010011, 32'b0000000??????????001?????0111011, 32'b000000???????????001?????0011011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_SLL_1;
      end
      32'b0000000??????????101?????0110011, 32'b000000???????????101?????0010011, 32'b0000000??????????101?????0111011, 32'b000000???????????101?????0011011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_SRL_1;
      end
      32'b0100000??????????101?????0110011, 32'b010000???????????101?????0010011, 32'b0100000??????????101?????0111011, 32'b010000???????????101?????0011011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_SRA_1;
      end
      32'b0000000??????????111?????0110011, 32'b?????????????????111?????0010011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_AND_1;
      end
      32'b0000000??????????110?????0110011, 32'b?????????????????110?????0010011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_OR_1;
      end
      32'b?????????????????????????0110111 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_LUI;
      end
      32'b?????????????????????????0010111 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_AUIPC;
      end
      32'b??????????0??????????????1101111 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_JAL;
      end
      32'b?????????????????000?????1100111 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_JALR;
      end
      32'b?????????????????000???0?1100011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_BEQ;
      end
      32'b?????????????????001???0?1100011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_BNE;
      end
      32'b?????????????????100???0?1100011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_BLT;
      end
      32'b?????????????????101???0?1100011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_BGE;
      end
      32'b?????????????????110???0?1100011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_BLTU;
      end
      32'b?????????????????111???0?1100011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_BGEU;
      end
      32'b?????????????????001?????1110011, 32'b?????????????????010?????1110011, 32'b?????????????????011?????1110011, 32'b?????????????????101?????1110011, 32'b?????????????????110?????1110011, 32'b?????????????????111?????1110011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_CSR;
      end
      default : begin
        decode_DecodePlugin_alu_ctrl = 5'h0;
      end
    endcase
  end

  always @(*) begin
    casez(decode_INSTRUCTION)
      32'b?????????????????000?????0000011 : begin
        decode_DecodePlugin_mem_ctrl = MemCtrlEnum_LB;
      end
      32'b?????????????????100?????0000011 : begin
        decode_DecodePlugin_mem_ctrl = MemCtrlEnum_LBU;
      end
      32'b?????????????????001?????0000011 : begin
        decode_DecodePlugin_mem_ctrl = MemCtrlEnum_LH;
      end
      32'b?????????????????101?????0000011 : begin
        decode_DecodePlugin_mem_ctrl = MemCtrlEnum_LHU;
      end
      32'b?????????????????010?????0000011 : begin
        decode_DecodePlugin_mem_ctrl = MemCtrlEnum_LW;
      end
      32'b?????????????????110?????0000011 : begin
        decode_DecodePlugin_mem_ctrl = MemCtrlEnum_LWU;
      end
      32'b?????????????????011?????0000011 : begin
        decode_DecodePlugin_mem_ctrl = MemCtrlEnum_LD;
      end
      32'b?????????????????000?????0100011 : begin
        decode_DecodePlugin_mem_ctrl = MemCtrlEnum_SB;
      end
      32'b?????????????????001?????0100011 : begin
        decode_DecodePlugin_mem_ctrl = MemCtrlEnum_SH;
      end
      32'b?????????????????010?????0100011 : begin
        decode_DecodePlugin_mem_ctrl = MemCtrlEnum_SW;
      end
      32'b?????????????????011?????0100011 : begin
        decode_DecodePlugin_mem_ctrl = MemCtrlEnum_SD;
      end
      default : begin
        decode_DecodePlugin_mem_ctrl = 4'b0000;
      end
    endcase
  end

  always @(*) begin
    casez(decode_INSTRUCTION)
      32'b?????????????????000?????0000011 : begin
        decode_DecodePlugin_is_load = 1'b1;
      end
      32'b?????????????????100?????0000011 : begin
        decode_DecodePlugin_is_load = 1'b1;
      end
      32'b?????????????????001?????0000011 : begin
        decode_DecodePlugin_is_load = 1'b1;
      end
      32'b?????????????????101?????0000011 : begin
        decode_DecodePlugin_is_load = 1'b1;
      end
      32'b?????????????????010?????0000011 : begin
        decode_DecodePlugin_is_load = 1'b1;
      end
      32'b?????????????????110?????0000011 : begin
        decode_DecodePlugin_is_load = 1'b1;
      end
      32'b?????????????????011?????0000011 : begin
        decode_DecodePlugin_is_load = 1'b1;
      end
      32'b?????????????????000?????0100011 : begin
        decode_DecodePlugin_is_load = 1'b0;
      end
      32'b?????????????????001?????0100011 : begin
        decode_DecodePlugin_is_load = 1'b0;
      end
      32'b?????????????????010?????0100011 : begin
        decode_DecodePlugin_is_load = 1'b0;
      end
      32'b?????????????????011?????0100011 : begin
        decode_DecodePlugin_is_load = 1'b0;
      end
      default : begin
        decode_DecodePlugin_is_load = 1'b0;
      end
    endcase
  end

  always @(*) begin
    casez(decode_INSTRUCTION)
      32'b?????????????????000?????0000011 : begin
        decode_DecodePlugin_is_store = 1'b0;
      end
      32'b?????????????????100?????0000011 : begin
        decode_DecodePlugin_is_store = 1'b0;
      end
      32'b?????????????????001?????0000011 : begin
        decode_DecodePlugin_is_store = 1'b0;
      end
      32'b?????????????????101?????0000011 : begin
        decode_DecodePlugin_is_store = 1'b0;
      end
      32'b?????????????????010?????0000011 : begin
        decode_DecodePlugin_is_store = 1'b0;
      end
      32'b?????????????????110?????0000011 : begin
        decode_DecodePlugin_is_store = 1'b0;
      end
      32'b?????????????????011?????0000011 : begin
        decode_DecodePlugin_is_store = 1'b0;
      end
      32'b?????????????????000?????0100011 : begin
        decode_DecodePlugin_is_store = 1'b1;
      end
      32'b?????????????????001?????0100011 : begin
        decode_DecodePlugin_is_store = 1'b1;
      end
      32'b?????????????????010?????0100011 : begin
        decode_DecodePlugin_is_store = 1'b1;
      end
      32'b?????????????????011?????0100011 : begin
        decode_DecodePlugin_is_store = 1'b1;
      end
      default : begin
        decode_DecodePlugin_is_store = 1'b0;
      end
    endcase
  end

  always @(*) begin
    casez(decode_INSTRUCTION)
      32'b00000000000000000000000001110011 : begin
        decode_DecodePlugin_csr_ctrl = CsrCtrlEnum_ECALL;
      end
      32'b00000000000100000000000001110011 : begin
        decode_DecodePlugin_csr_ctrl = CsrCtrlEnum_EBREAK;
      end
      32'b00110000001000000000000001110011 : begin
        decode_DecodePlugin_csr_ctrl = CsrCtrlEnum_MRET;
      end
      32'b?????????????????001?????1110011 : begin
        decode_DecodePlugin_csr_ctrl = CsrCtrlEnum_CSRRW;
      end
      32'b?????????????????010?????1110011 : begin
        decode_DecodePlugin_csr_ctrl = CsrCtrlEnum_CSRRS;
      end
      32'b?????????????????011?????1110011 : begin
        decode_DecodePlugin_csr_ctrl = CsrCtrlEnum_CSRRC;
      end
      32'b?????????????????101?????1110011 : begin
        decode_DecodePlugin_csr_ctrl = CsrCtrlEnum_CSRRWI;
      end
      32'b?????????????????110?????1110011 : begin
        decode_DecodePlugin_csr_ctrl = CsrCtrlEnum_CSRRSI;
      end
      32'b?????????????????111?????1110011 : begin
        decode_DecodePlugin_csr_ctrl = CsrCtrlEnum_CSRRCI;
      end
      default : begin
        decode_DecodePlugin_csr_ctrl = 4'b0000;
      end
    endcase
  end

  assign decode_DecodePlugin_rs1 = regFileModule_1_read_ports_rs1_value;
  assign decode_DecodePlugin_rs2 = regFileModule_1_read_ports_rs2_value;
  assign decode_DecodePlugin_rd_wen = ((((((! (decode_INSTRUCTION[6 : 0] == 7'h23)) && (! (decode_INSTRUCTION[6 : 0] == 7'h63))) && (! ((decode_INSTRUCTION & 32'hffffffff) == 32'h00100073))) && (! ((decode_INSTRUCTION & 32'hffffffff) == 32'h00000073))) && (! ((decode_INSTRUCTION & 32'hffffffff) == 32'h30200073))) && (decode_INSTRUCTION[6 : 0] != 7'h0f));
  assign DecodePlugin_hazard_decode_rs1_req = decode_DecodePlugin_rs1_req;
  assign DecodePlugin_hazard_decode_rs2_req = decode_DecodePlugin_rs2_req;
  assign DecodePlugin_hazard_decode_rs1_addr = decode_DecodePlugin_rs1_addr;
  assign DecodePlugin_hazard_decode_rs2_addr = decode_DecodePlugin_rs2_addr;
  assign regFileModule_1_write_ports_rd_wen = (writeback_arbitration_isFiring && _zz_DecodePlugin_hazard_rs1_from_wb_1);
  assign execute_ALUPlugin_src1_word = execute_ALUPlugin_src1[31 : 0];
  assign execute_ALUPlugin_src2_word = execute_ALUPlugin_src2[31 : 0];
  assign execute_ALUPlugin_shift_bits = execute_ALUPlugin_src2[5 : 0];
  assign execute_ALUPlugin_add_result = ($signed(_zz_execute_ALUPlugin_add_result) + $signed(_zz_execute_ALUPlugin_add_result_1));
  assign execute_ALUPlugin_sub_result = ($signed(_zz_execute_ALUPlugin_sub_result) - $signed(_zz_execute_ALUPlugin_sub_result_1));
  assign execute_ALUPlugin_slt_result = ($signed(_zz_execute_ALUPlugin_slt_result) < $signed(_zz_execute_ALUPlugin_slt_result_1));
  assign execute_ALUPlugin_sltu_result = (execute_ALUPlugin_src1 < execute_ALUPlugin_src2);
  assign execute_ALUPlugin_xor_result = (execute_ALUPlugin_src1 ^ execute_ALUPlugin_src2);
  assign execute_ALUPlugin_sll_result = (execute_ALUPlugin_src1 <<< execute_ALUPlugin_shift_bits);
  assign execute_ALUPlugin_srl_result = (execute_ALUPlugin_src1 >>> execute_ALUPlugin_shift_bits);
  assign execute_ALUPlugin_sra_result = ($signed(_zz_execute_ALUPlugin_sra_result) >>> execute_ALUPlugin_shift_bits);
  assign execute_ALUPlugin_and_result = (execute_ALUPlugin_src1 & execute_ALUPlugin_src2);
  assign execute_ALUPlugin_or_result = (execute_ALUPlugin_src1 | execute_ALUPlugin_src2);
  assign _zz_execute_ALUPlugin_addw_result = execute_ALUPlugin_add_result[31];
  always @(*) begin
    _zz_execute_ALUPlugin_addw_result_1[31] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[30] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[29] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[28] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[27] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[26] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[25] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[24] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[23] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[22] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[21] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[20] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[19] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[18] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[17] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[16] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[15] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[14] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[13] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[12] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[11] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[10] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[9] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[8] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[7] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[6] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[5] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[4] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[3] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[2] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[1] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[0] = _zz_execute_ALUPlugin_addw_result;
  end

  assign execute_ALUPlugin_addw_result = {_zz_execute_ALUPlugin_addw_result_1,_zz_execute_ALUPlugin_addw_result_2};
  assign _zz_execute_ALUPlugin_subw_result = execute_ALUPlugin_sub_result[31];
  always @(*) begin
    _zz_execute_ALUPlugin_subw_result_1[31] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[30] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[29] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[28] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[27] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[26] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[25] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[24] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[23] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[22] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[21] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[20] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[19] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[18] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[17] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[16] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[15] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[14] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[13] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[12] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[11] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[10] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[9] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[8] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[7] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[6] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[5] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[4] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[3] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[2] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[1] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[0] = _zz_execute_ALUPlugin_subw_result;
  end

  assign execute_ALUPlugin_subw_result = {_zz_execute_ALUPlugin_subw_result_1,_zz_execute_ALUPlugin_subw_result_2};
  assign execute_ALUPlugin_sllw_temp = (execute_ALUPlugin_src1_word <<< execute_ALUPlugin_shift_bits[4 : 0]);
  assign _zz_execute_ALUPlugin_sllw_result = execute_ALUPlugin_sllw_temp[31];
  always @(*) begin
    _zz_execute_ALUPlugin_sllw_result_1[31] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[30] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[29] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[28] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[27] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[26] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[25] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[24] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[23] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[22] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[21] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[20] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[19] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[18] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[17] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[16] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[15] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[14] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[13] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[12] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[11] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[10] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[9] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[8] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[7] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[6] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[5] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[4] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[3] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[2] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[1] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[0] = _zz_execute_ALUPlugin_sllw_result;
  end

  assign execute_ALUPlugin_sllw_result = {_zz_execute_ALUPlugin_sllw_result_1,execute_ALUPlugin_sllw_temp};
  assign execute_ALUPlugin_srlw_temp = (execute_ALUPlugin_src1_word >>> execute_ALUPlugin_shift_bits[4 : 0]);
  assign _zz_execute_ALUPlugin_srlw_result = execute_ALUPlugin_srlw_temp[31];
  always @(*) begin
    _zz_execute_ALUPlugin_srlw_result_1[31] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[30] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[29] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[28] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[27] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[26] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[25] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[24] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[23] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[22] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[21] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[20] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[19] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[18] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[17] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[16] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[15] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[14] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[13] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[12] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[11] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[10] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[9] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[8] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[7] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[6] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[5] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[4] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[3] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[2] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[1] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[0] = _zz_execute_ALUPlugin_srlw_result;
  end

  assign execute_ALUPlugin_srlw_result = {_zz_execute_ALUPlugin_srlw_result_1,execute_ALUPlugin_srlw_temp};
  assign execute_ALUPlugin_sraw_temp = ($signed(_zz_execute_ALUPlugin_sraw_temp) >>> execute_ALUPlugin_shift_bits[4 : 0]);
  assign _zz_execute_ALUPlugin_sraw_result = execute_ALUPlugin_sraw_temp[31];
  always @(*) begin
    _zz_execute_ALUPlugin_sraw_result_1[31] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[30] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[29] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[28] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[27] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[26] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[25] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[24] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[23] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[22] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[21] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[20] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[19] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[18] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[17] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[16] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[15] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[14] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[13] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[12] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[11] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[10] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[9] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[8] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[7] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[6] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[5] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[4] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[3] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[2] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[1] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[0] = _zz_execute_ALUPlugin_sraw_result;
  end

  assign execute_ALUPlugin_sraw_result = {_zz_execute_ALUPlugin_sraw_result_1,execute_ALUPlugin_sraw_temp};
  assign execute_ALUPlugin_jal = (execute_ALU_CTRL == AluCtrlEnum_JAL);
  assign execute_ALUPlugin_jalr = (execute_ALU_CTRL == AluCtrlEnum_JALR);
  assign execute_ALUPlugin_beq = (execute_ALU_CTRL == AluCtrlEnum_BEQ);
  assign execute_ALUPlugin_bne = (execute_ALU_CTRL == AluCtrlEnum_BNE);
  assign execute_ALUPlugin_blt = (execute_ALU_CTRL == AluCtrlEnum_BLT);
  assign execute_ALUPlugin_bge = (execute_ALU_CTRL == AluCtrlEnum_BGE);
  assign execute_ALUPlugin_bltu = (execute_ALU_CTRL == AluCtrlEnum_BLTU);
  assign execute_ALUPlugin_bgeu = (execute_ALU_CTRL == AluCtrlEnum_BGEU);
  assign execute_ALUPlugin_branch_or_jalr = ((((((execute_ALUPlugin_jalr || execute_ALUPlugin_beq) || execute_ALUPlugin_bne) || execute_ALUPlugin_blt) || execute_ALUPlugin_bge) || execute_ALUPlugin_bltu) || execute_ALUPlugin_bgeu);
  assign execute_ALUPlugin_branch_or_jump = (execute_ALUPlugin_branch_or_jalr || execute_ALUPlugin_jal);
  assign execute_ALUPlugin_rd_is_link = ((execute_RD_ADDR == 5'h0) || (execute_RD_ADDR == 5'h05));
  assign execute_ALUPlugin_rs1_is_link = ((execute_RS1_ADDR == 5'h0) || (execute_RS1_ADDR == 5'h05));
  always @(*) begin
    execute_ALUPlugin_is_call = 1'b0;
    if(execute_ALUPlugin_jal) begin
      if(execute_ALUPlugin_rd_is_link) begin
        execute_ALUPlugin_is_call = 1'b1;
      end else begin
        execute_ALUPlugin_is_call = 1'b0;
      end
    end else begin
      if(execute_ALUPlugin_jalr) begin
        if(execute_ALUPlugin_rd_is_link) begin
          if(execute_ALUPlugin_rs1_is_link) begin
            if(when_AluPlugin_l270) begin
              execute_ALUPlugin_is_call = 1'b1;
            end else begin
              execute_ALUPlugin_is_call = 1'b1;
            end
          end else begin
            execute_ALUPlugin_is_call = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    execute_ALUPlugin_is_ret = 1'b0;
    if(execute_ALUPlugin_jal) begin
      if(execute_ALUPlugin_rd_is_link) begin
        execute_ALUPlugin_is_ret = 1'b0;
      end else begin
        execute_ALUPlugin_is_ret = 1'b0;
      end
    end else begin
      if(execute_ALUPlugin_jalr) begin
        if(execute_ALUPlugin_rd_is_link) begin
          if(execute_ALUPlugin_rs1_is_link) begin
            if(!when_AluPlugin_l270) begin
              execute_ALUPlugin_is_ret = 1'b1;
            end
          end
        end else begin
          if(execute_ALUPlugin_rs1_is_link) begin
            execute_ALUPlugin_is_ret = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    execute_ALUPlugin_is_jmp = 1'b0;
    if(execute_ALUPlugin_jal) begin
      if(execute_ALUPlugin_rd_is_link) begin
        execute_ALUPlugin_is_jmp = 1'b0;
      end else begin
        execute_ALUPlugin_is_jmp = 1'b1;
      end
    end else begin
      if(execute_ALUPlugin_jalr) begin
        if(!execute_ALUPlugin_rd_is_link) begin
          if(!execute_ALUPlugin_rs1_is_link) begin
            execute_ALUPlugin_is_jmp = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    execute_ALUPlugin_redirect_pc_next = (execute_PC + 64'h0000000000000004);
    if(execute_ALUPlugin_branch_or_jump) begin
      if(execute_ALUPlugin_branch_taken) begin
        if(when_AluPlugin_l234) begin
          execute_ALUPlugin_redirect_pc_next = execute_ALUPlugin_pc_next;
        end
      end else begin
        if(execute_PREDICT_TAKEN) begin
          execute_ALUPlugin_redirect_pc_next = (execute_PC + 64'h0000000000000004);
        end
      end
    end
  end

  always @(*) begin
    execute_ALUPlugin_redirect_valid = 1'b0;
    if(execute_ALUPlugin_branch_or_jump) begin
      if(execute_ALUPlugin_branch_taken) begin
        if(when_AluPlugin_l234) begin
          execute_ALUPlugin_redirect_valid = execute_arbitration_isFiring;
        end
      end else begin
        if(execute_PREDICT_TAKEN) begin
          execute_ALUPlugin_redirect_valid = execute_arbitration_isFiring;
        end
      end
    end
  end

  assign when_AluPlugin_l77 = (((execute_ALU_CTRL == AluCtrlEnum_AUIPC) || execute_ALUPlugin_jal) || execute_ALUPlugin_jalr);
  always @(*) begin
    if(when_AluPlugin_l77) begin
      execute_ALUPlugin_src1 = execute_PC;
    end else begin
      if(execute_RS1_FROM_MEM) begin
        execute_ALUPlugin_src1 = memaccess_ALU_RESULT;
      end else begin
        if(execute_RS1_FROM_LOAD) begin
          execute_ALUPlugin_src1 = memaccess_LSU_RDATA;
        end else begin
          if(execute_RS1_FROM_WB) begin
            execute_ALUPlugin_src1 = _zz_execute_MEM_WDATA_2;
          end else begin
            execute_ALUPlugin_src1 = execute_RS1;
          end
        end
      end
    end
  end

  assign when_AluPlugin_l95 = (execute_ALUPlugin_jal || execute_ALUPlugin_jalr);
  always @(*) begin
    if(when_AluPlugin_l95) begin
      execute_ALUPlugin_src2 = 64'h0000000000000004;
    end else begin
      if(execute_SRC2_IS_IMM) begin
        execute_ALUPlugin_src2 = execute_IMM;
      end else begin
        if(execute_RS2_FROM_MEM) begin
          execute_ALUPlugin_src2 = memaccess_ALU_RESULT;
        end else begin
          if(execute_RS2_FROM_LOAD) begin
            execute_ALUPlugin_src2 = memaccess_LSU_RDATA;
          end else begin
            if(execute_RS2_FROM_WB) begin
              execute_ALUPlugin_src2 = _zz_execute_MEM_WDATA_2;
            end else begin
              execute_ALUPlugin_src2 = execute_RS2;
            end
          end
        end
      end
    end
  end

  always @(*) begin
    if(execute_CTRL_RS1_FROM_MEM) begin
      execute_ALUPlugin_branch_src1 = _zz_execute_MEM_WDATA_1;
    end else begin
      if(execute_CTRL_RS1_FROM_LOAD) begin
        execute_ALUPlugin_branch_src1 = _zz_execute_MEM_WDATA;
      end else begin
        if(execute_CTRL_RS1_FROM_WB) begin
          execute_ALUPlugin_branch_src1 = _zz_execute_MEM_WDATA_2;
        end else begin
          execute_ALUPlugin_branch_src1 = execute_RS1;
        end
      end
    end
  end

  always @(*) begin
    if(execute_CTRL_RS2_FROM_MEM) begin
      execute_ALUPlugin_branch_src2 = _zz_execute_MEM_WDATA_1;
    end else begin
      if(execute_CTRL_RS2_FROM_LOAD) begin
        execute_ALUPlugin_branch_src2 = _zz_execute_MEM_WDATA;
      end else begin
        if(execute_CTRL_RS2_FROM_WB) begin
          execute_ALUPlugin_branch_src2 = _zz_execute_MEM_WDATA_2;
        end else begin
          execute_ALUPlugin_branch_src2 = execute_RS2;
        end
      end
    end
  end

  assign when_AluPlugin_l146 = (execute_ALU_WORD == 1'b1);
  always @(*) begin
    if((execute_ALU_CTRL == AluCtrlEnum_ADD)) begin
        if(when_AluPlugin_l146) begin
          execute_ALUPlugin_alu_result = execute_ALUPlugin_addw_result;
        end else begin
          execute_ALUPlugin_alu_result = execute_ALUPlugin_add_result;
        end
    end else if((execute_ALU_CTRL == AluCtrlEnum_SUB)) begin
        if(when_AluPlugin_l153) begin
          execute_ALUPlugin_alu_result = execute_ALUPlugin_subw_result;
        end else begin
          execute_ALUPlugin_alu_result = execute_ALUPlugin_sub_result;
        end
    end else if((execute_ALU_CTRL == AluCtrlEnum_SLT)) begin
        execute_ALUPlugin_alu_result = {_zz_execute_ALUPlugin_alu_result,execute_ALUPlugin_slt_result};
    end else if((execute_ALU_CTRL == AluCtrlEnum_SLTU)) begin
        execute_ALUPlugin_alu_result = {_zz_execute_ALUPlugin_alu_result_1,execute_ALUPlugin_sltu_result};
    end else if((execute_ALU_CTRL == AluCtrlEnum_XOR_1)) begin
        execute_ALUPlugin_alu_result = execute_ALUPlugin_xor_result;
    end else if((execute_ALU_CTRL == AluCtrlEnum_SLL_1)) begin
        if(when_AluPlugin_l169) begin
          execute_ALUPlugin_alu_result = execute_ALUPlugin_sllw_result;
        end else begin
          execute_ALUPlugin_alu_result = execute_ALUPlugin_sll_result;
        end
    end else if((execute_ALU_CTRL == AluCtrlEnum_SRL_1)) begin
        if(when_AluPlugin_l176) begin
          execute_ALUPlugin_alu_result = execute_ALUPlugin_srlw_result;
        end else begin
          execute_ALUPlugin_alu_result = execute_ALUPlugin_srl_result;
        end
    end else if((execute_ALU_CTRL == AluCtrlEnum_SRA_1)) begin
        if(when_AluPlugin_l183) begin
          execute_ALUPlugin_alu_result = execute_ALUPlugin_sraw_result;
        end else begin
          execute_ALUPlugin_alu_result = execute_ALUPlugin_sra_result;
        end
    end else if((execute_ALU_CTRL == AluCtrlEnum_AND_1)) begin
        execute_ALUPlugin_alu_result = execute_ALUPlugin_and_result;
    end else if((execute_ALU_CTRL == AluCtrlEnum_OR_1)) begin
        execute_ALUPlugin_alu_result = execute_ALUPlugin_or_result;
    end else if((execute_ALU_CTRL == AluCtrlEnum_LUI)) begin
        execute_ALUPlugin_alu_result = execute_IMM;
    end else if((execute_ALU_CTRL == AluCtrlEnum_JAL) || (execute_ALU_CTRL == AluCtrlEnum_JALR) || (execute_ALU_CTRL == AluCtrlEnum_AUIPC)) begin
        execute_ALUPlugin_alu_result = execute_ALUPlugin_add_result;
    end else if((execute_ALU_CTRL == AluCtrlEnum_CSR)) begin
        execute_ALUPlugin_alu_result = execute_CSR_RDATA;
    end else begin
        execute_ALUPlugin_alu_result = execute_ALUPlugin_add_result;
    end
  end

  assign when_AluPlugin_l153 = (execute_ALU_WORD == 1'b1);
  assign _zz_execute_ALUPlugin_alu_result[62 : 0] = 63'h0;
  assign _zz_execute_ALUPlugin_alu_result_1[62 : 0] = 63'h0;
  assign when_AluPlugin_l169 = (execute_ALU_WORD == 1'b1);
  assign when_AluPlugin_l176 = (execute_ALU_WORD == 1'b1);
  assign when_AluPlugin_l183 = (execute_ALU_WORD == 1'b1);
  assign execute_ALUPlugin_beq_result = (execute_ALUPlugin_beq && (execute_ALUPlugin_branch_src1 == execute_ALUPlugin_branch_src2));
  assign execute_ALUPlugin_bne_result = (execute_ALUPlugin_bne && (execute_ALUPlugin_branch_src1 != execute_ALUPlugin_branch_src2));
  assign execute_ALUPlugin_blt_result = (execute_ALUPlugin_blt && ($signed(_zz_execute_ALUPlugin_blt_result) < $signed(_zz_execute_ALUPlugin_blt_result_1)));
  assign execute_ALUPlugin_bge_result = (execute_ALUPlugin_bge && ($signed(_zz_execute_ALUPlugin_bge_result) <= $signed(_zz_execute_ALUPlugin_bge_result_1)));
  assign execute_ALUPlugin_bltu_result = (execute_ALUPlugin_bltu && (execute_ALUPlugin_branch_src1 < execute_ALUPlugin_branch_src2));
  assign execute_ALUPlugin_bgeu_result = (execute_ALUPlugin_bgeu && (execute_ALUPlugin_branch_src2 <= execute_ALUPlugin_branch_src1));
  assign execute_ALUPlugin_branch_taken = (((((((execute_ALUPlugin_beq_result || execute_ALUPlugin_bne_result) || execute_ALUPlugin_blt_result) || execute_ALUPlugin_bge_result) || execute_ALUPlugin_bltu_result) || execute_ALUPlugin_bgeu_result) || execute_ALUPlugin_jal) || execute_ALUPlugin_jalr);
  assign when_AluPlugin_l226 = (execute_ALU_CTRL == AluCtrlEnum_JALR);
  always @(*) begin
    if(when_AluPlugin_l226) begin
      execute_ALUPlugin_pc_next = _zz_execute_ALUPlugin_pc_next;
    end else begin
      execute_ALUPlugin_pc_next = _zz_execute_ALUPlugin_pc_next_6;
    end
  end

  assign when_AluPlugin_l234 = ((! execute_PREDICT_TAKEN) || (execute_PC_NEXT != execute_ALUPlugin_pc_next));
  assign when_AluPlugin_l270 = (execute_RD_ADDR == execute_RS1_ADDR);
  assign DecodePlugin_hazard_rs1_from_mem = ((((memaccess_arbitration_isValid && _zz_DecodePlugin_hazard_rs1_from_mem_3) && (_zz_DecodePlugin_hazard_rs1_from_mem_2 != 5'h0)) && (_zz_DecodePlugin_hazard_rs1_from_mem_2 == _zz_DecodePlugin_hazard_rs1_from_mem_1)) && (! _zz_DecodePlugin_hazard_rs1_from_mem));
  assign DecodePlugin_hazard_rs2_from_mem = ((((memaccess_arbitration_isValid && _zz_DecodePlugin_hazard_rs1_from_mem_3) && (_zz_DecodePlugin_hazard_rs1_from_mem_2 != 5'h0)) && (_zz_DecodePlugin_hazard_rs1_from_mem_2 == _zz_DecodePlugin_hazard_rs2_from_mem)) && (! _zz_DecodePlugin_hazard_rs1_from_mem));
  assign DecodePlugin_hazard_rs1_from_load = ((((memaccess_arbitration_isValid && _zz_DecodePlugin_hazard_rs1_from_mem_3) && (_zz_DecodePlugin_hazard_rs1_from_mem_2 != 5'h0)) && (_zz_DecodePlugin_hazard_rs1_from_mem_2 == _zz_DecodePlugin_hazard_rs1_from_mem_1)) && _zz_DecodePlugin_hazard_rs1_from_mem);
  assign DecodePlugin_hazard_rs2_from_load = ((((memaccess_arbitration_isValid && _zz_DecodePlugin_hazard_rs1_from_mem_3) && (_zz_DecodePlugin_hazard_rs1_from_mem_2 != 5'h0)) && (_zz_DecodePlugin_hazard_rs1_from_mem_2 == _zz_DecodePlugin_hazard_rs2_from_mem)) && _zz_DecodePlugin_hazard_rs1_from_mem);
  assign DecodePlugin_hazard_rs1_from_wb = ((((writeback_arbitration_isValid && _zz_DecodePlugin_hazard_rs1_from_wb_1) && (_zz_DecodePlugin_hazard_rs1_from_wb != 5'h0)) && (_zz_DecodePlugin_hazard_rs1_from_wb == _zz_DecodePlugin_hazard_rs1_from_mem_1)) && (! (DecodePlugin_hazard_rs1_from_mem || DecodePlugin_hazard_rs1_from_load)));
  assign DecodePlugin_hazard_rs2_from_wb = ((((writeback_arbitration_isValid && _zz_DecodePlugin_hazard_rs1_from_wb_1) && (_zz_DecodePlugin_hazard_rs1_from_wb != 5'h0)) && (_zz_DecodePlugin_hazard_rs1_from_wb == _zz_DecodePlugin_hazard_rs2_from_mem)) && (! (DecodePlugin_hazard_rs2_from_mem || DecodePlugin_hazard_rs2_from_load)));
  assign DecodePlugin_hazard_load_use = ((memaccess_arbitration_isValid && _zz_DecodePlugin_hazard_rs1_from_mem) && (((_zz_DecodePlugin_hazard_rs1_from_mem_2 == _zz_DecodePlugin_hazard_rs1_from_mem_1) && (! DecodePlugin_hazard_rs1_from_wb)) || ((_zz_DecodePlugin_hazard_rs1_from_mem_2 == _zz_DecodePlugin_hazard_rs2_from_mem) && (! DecodePlugin_hazard_rs2_from_wb))));
  assign DecodePlugin_hazard_ctrl_rs1_from_mem = ((execute_arbitration_isValid && _zz_DecodePlugin_hazard_ctrl_rs1_from_mem) && DecodePlugin_hazard_rs1_from_mem);
  assign DecodePlugin_hazard_ctrl_rs2_from_mem = ((execute_arbitration_isValid && _zz_DecodePlugin_hazard_ctrl_rs1_from_mem) && DecodePlugin_hazard_rs2_from_mem);
  assign DecodePlugin_hazard_ctrl_rs1_from_load = ((execute_arbitration_isValid && _zz_DecodePlugin_hazard_ctrl_rs1_from_mem) && DecodePlugin_hazard_rs1_from_load);
  assign DecodePlugin_hazard_ctrl_rs2_from_load = ((execute_arbitration_isValid && _zz_DecodePlugin_hazard_ctrl_rs1_from_mem) && DecodePlugin_hazard_rs2_from_load);
  assign DecodePlugin_hazard_ctrl_rs1_from_wb = ((execute_arbitration_isValid && _zz_DecodePlugin_hazard_ctrl_rs1_from_mem) && DecodePlugin_hazard_rs1_from_wb);
  assign DecodePlugin_hazard_ctrl_rs2_from_wb = ((execute_arbitration_isValid && _zz_DecodePlugin_hazard_ctrl_rs1_from_mem) && DecodePlugin_hazard_rs2_from_wb);
  assign DecodePlugin_hazard_ctrl_load_use = ((execute_arbitration_isValid && _zz_DecodePlugin_hazard_ctrl_rs1_from_mem) && DecodePlugin_hazard_load_use);
  assign fetch_arbitration_haltItself = 1'b0;
  assign fetch_arbitration_flushIt = (when_FetchPlugin_l97 || when_FetchPlugin_l94);
  assign decode_arbitration_haltItself = 1'b0;
  assign decode_arbitration_flushIt = (when_FetchPlugin_l97 || when_FetchPlugin_l94);
  assign execute_arbitration_haltItself = execute_INT_HOLD;
  assign execute_arbitration_flushIt = 1'b0;
  assign memaccess_arbitration_haltItself = _zz_memaccess_arbitration_haltItself;
  assign memaccess_arbitration_flushIt = 1'b0;
  assign writeback_arbitration_haltItself = _zz_memaccess_arbitration_haltItself;
  assign writeback_arbitration_flushIt = 1'b0;
  assign clint_1_ecall = (execute_arbitration_isValid && (_zz_ecall == CsrCtrlEnum_ECALL));
  assign clint_1_ebreak = (execute_arbitration_isValid && (_zz_ecall == CsrCtrlEnum_EBREAK));
  assign clint_1_mret = (execute_arbitration_isValid && (_zz_ecall == CsrCtrlEnum_MRET));
  assign execute_ExcepPlugin_csrrs_wdata = (execute_SRC1 | execute_CSR_RDATA);
  assign execute_ExcepPlugin_csrrc_wdata = ((~ execute_SRC1) & execute_CSR_RDATA);
  assign execute_ExcepPlugin_csrrsi_wdata = (execute_IMM | execute_CSR_RDATA);
  assign execute_ExcepPlugin_csrrci_wdata = ((~ execute_IMM) & execute_CSR_RDATA);
  always @(*) begin
    if((execute_CSR_CTRL == CsrCtrlEnum_CSRRW)) begin
        execute_ExcepPlugin_csr_wdata = execute_SRC1;
    end else if((execute_CSR_CTRL == CsrCtrlEnum_CSRRS)) begin
        execute_ExcepPlugin_csr_wdata = execute_ExcepPlugin_csrrs_wdata;
    end else if((execute_CSR_CTRL == CsrCtrlEnum_CSRRC)) begin
        execute_ExcepPlugin_csr_wdata = execute_ExcepPlugin_csrrc_wdata;
    end else if((execute_CSR_CTRL == CsrCtrlEnum_CSRRWI)) begin
        execute_ExcepPlugin_csr_wdata = execute_IMM;
    end else if((execute_CSR_CTRL == CsrCtrlEnum_CSRRSI)) begin
        execute_ExcepPlugin_csr_wdata = execute_ExcepPlugin_csrrsi_wdata;
    end else if((execute_CSR_CTRL == CsrCtrlEnum_CSRRCI)) begin
        execute_ExcepPlugin_csr_wdata = execute_ExcepPlugin_csrrci_wdata;
    end else begin
        execute_ExcepPlugin_csr_wdata = 64'h0;
    end
  end

  assign timer_1_addr = _zz_execute_MEM_WDATA_1;
  assign memaccess_LSUPlugin_cpu_addr = memaccess_ALU_RESULT;
  assign memaccess_LSUPlugin_cpu_addr_offset = memaccess_LSUPlugin_cpu_addr[2 : 0];
  assign memaccess_LSUPlugin_is_mem = (memaccess_IS_LOAD || memaccess_IS_STORE);
  assign memaccess_LSUPlugin_is_timer = ((memaccess_LSUPlugin_cpu_addr == 64'h000000000200bff8) || (memaccess_LSUPlugin_cpu_addr == 64'h0000000002004000));
  assign memaccess_LSUPlugin_dcache_rdata = (DCachePlugin_dcache_access_rsp_payload_data >>> _zz_memaccess_LSUPlugin_dcache_rdata);
  assign _zz_memaccess_LSUPlugin_dcache_lb = memaccess_LSUPlugin_dcache_rdata[7];
  always @(*) begin
    _zz_memaccess_LSUPlugin_dcache_lb_1[55] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[54] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[53] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[52] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[51] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[50] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[49] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[48] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[47] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[46] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[45] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[44] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[43] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[42] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[41] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[40] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[39] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[38] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[37] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[36] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[35] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[34] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[33] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[32] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[31] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[30] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[29] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[28] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[27] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[26] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[25] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[24] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[23] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[22] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[21] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[20] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[19] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[18] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[17] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[16] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[15] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[14] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[13] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[12] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[11] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[10] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[9] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[8] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[7] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[6] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[5] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[4] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[3] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[2] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[1] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[0] = _zz_memaccess_LSUPlugin_dcache_lb;
  end

  assign memaccess_LSUPlugin_dcache_lb = {_zz_memaccess_LSUPlugin_dcache_lb_1,memaccess_LSUPlugin_dcache_rdata[7 : 0]};
  assign _zz_1 = zz__zz_memaccess_LSUPlugin_dcache_lbu(1'b0);
  always @(*) _zz_memaccess_LSUPlugin_dcache_lbu = _zz_1;
  assign memaccess_LSUPlugin_dcache_lbu = {_zz_memaccess_LSUPlugin_dcache_lbu,memaccess_LSUPlugin_dcache_rdata[7 : 0]};
  assign _zz_memaccess_LSUPlugin_dcache_lh = memaccess_LSUPlugin_dcache_rdata[15];
  always @(*) begin
    _zz_memaccess_LSUPlugin_dcache_lh_1[47] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[46] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[45] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[44] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[43] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[42] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[41] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[40] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[39] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[38] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[37] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[36] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[35] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[34] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[33] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[32] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[31] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[30] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[29] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[28] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[27] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[26] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[25] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[24] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[23] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[22] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[21] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[20] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[19] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[18] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[17] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[16] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[15] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[14] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[13] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[12] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[11] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[10] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[9] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[8] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[7] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[6] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[5] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[4] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[3] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[2] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[1] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[0] = _zz_memaccess_LSUPlugin_dcache_lh;
  end

  assign memaccess_LSUPlugin_dcache_lh = {_zz_memaccess_LSUPlugin_dcache_lh_1,memaccess_LSUPlugin_dcache_rdata[15 : 0]};
  assign _zz_2 = zz__zz_memaccess_LSUPlugin_dcache_lhu(1'b0);
  always @(*) _zz_memaccess_LSUPlugin_dcache_lhu = _zz_2;
  assign memaccess_LSUPlugin_dcache_lhu = {_zz_memaccess_LSUPlugin_dcache_lhu,memaccess_LSUPlugin_dcache_rdata[15 : 0]};
  assign _zz_memaccess_LSUPlugin_dcache_lw = memaccess_LSUPlugin_dcache_rdata[31];
  always @(*) begin
    _zz_memaccess_LSUPlugin_dcache_lw_1[31] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[30] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[29] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[28] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[27] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[26] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[25] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[24] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[23] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[22] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[21] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[20] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[19] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[18] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[17] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[16] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[15] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[14] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[13] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[12] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[11] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[10] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[9] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[8] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[7] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[6] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[5] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[4] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[3] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[2] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[1] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[0] = _zz_memaccess_LSUPlugin_dcache_lw;
  end

  assign memaccess_LSUPlugin_dcache_lw = {_zz_memaccess_LSUPlugin_dcache_lw_1,memaccess_LSUPlugin_dcache_rdata[31 : 0]};
  assign _zz_3 = zz__zz_memaccess_LSUPlugin_dcache_lwu(1'b0);
  always @(*) _zz_memaccess_LSUPlugin_dcache_lwu = _zz_3;
  assign memaccess_LSUPlugin_dcache_lwu = {_zz_memaccess_LSUPlugin_dcache_lwu,memaccess_LSUPlugin_dcache_rdata[31 : 0]};
  assign _zz_memaccess_LSUPlugin_dcache_sb = memaccess_MEM_WDATA[7];
  always @(*) begin
    _zz_memaccess_LSUPlugin_dcache_sb_1[55] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[54] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[53] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[52] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[51] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[50] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[49] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[48] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[47] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[46] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[45] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[44] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[43] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[42] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[41] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[40] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[39] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[38] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[37] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[36] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[35] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[34] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[33] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[32] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[31] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[30] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[29] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[28] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[27] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[26] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[25] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[24] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[23] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[22] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[21] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[20] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[19] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[18] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[17] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[16] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[15] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[14] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[13] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[12] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[11] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[10] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[9] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[8] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[7] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[6] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[5] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[4] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[3] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[2] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[1] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[0] = _zz_memaccess_LSUPlugin_dcache_sb;
  end

  assign memaccess_LSUPlugin_dcache_sb = {_zz_memaccess_LSUPlugin_dcache_sb_1,memaccess_MEM_WDATA[7 : 0]};
  assign _zz_memaccess_LSUPlugin_dcache_sh = memaccess_MEM_WDATA[15];
  always @(*) begin
    _zz_memaccess_LSUPlugin_dcache_sh_1[47] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[46] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[45] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[44] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[43] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[42] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[41] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[40] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[39] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[38] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[37] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[36] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[35] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[34] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[33] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[32] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[31] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[30] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[29] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[28] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[27] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[26] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[25] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[24] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[23] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[22] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[21] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[20] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[19] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[18] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[17] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[16] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[15] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[14] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[13] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[12] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[11] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[10] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[9] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[8] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[7] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[6] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[5] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[4] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[3] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[2] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[1] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[0] = _zz_memaccess_LSUPlugin_dcache_sh;
  end

  assign memaccess_LSUPlugin_dcache_sh = {_zz_memaccess_LSUPlugin_dcache_sh_1,memaccess_MEM_WDATA[15 : 0]};
  assign _zz_memaccess_LSUPlugin_dcache_sw = memaccess_MEM_WDATA[31];
  always @(*) begin
    _zz_memaccess_LSUPlugin_dcache_sw_1[31] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[30] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[29] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[28] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[27] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[26] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[25] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[24] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[23] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[22] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[21] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[20] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[19] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[18] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[17] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[16] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[15] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[14] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[13] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[12] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[11] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[10] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[9] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[8] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[7] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[6] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[5] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[4] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[3] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[2] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[1] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[0] = _zz_memaccess_LSUPlugin_dcache_sw;
  end

  assign memaccess_LSUPlugin_dcache_sw = {_zz_memaccess_LSUPlugin_dcache_sw_1,memaccess_MEM_WDATA[31 : 0]};
  assign memaccess_LSUPlugin_lsu_ready = 1'b1;
  always @(*) begin
    if((memaccess_MEM_CTRL == MemCtrlEnum_LB)) begin
        memaccess_LSUPlugin_dcache_data_load = memaccess_LSUPlugin_dcache_lb;
    end else if((memaccess_MEM_CTRL == MemCtrlEnum_LBU)) begin
        memaccess_LSUPlugin_dcache_data_load = memaccess_LSUPlugin_dcache_lbu;
    end else if((memaccess_MEM_CTRL == MemCtrlEnum_LH)) begin
        memaccess_LSUPlugin_dcache_data_load = memaccess_LSUPlugin_dcache_lh;
    end else if((memaccess_MEM_CTRL == MemCtrlEnum_LHU)) begin
        memaccess_LSUPlugin_dcache_data_load = memaccess_LSUPlugin_dcache_lhu;
    end else if((memaccess_MEM_CTRL == MemCtrlEnum_LW)) begin
        memaccess_LSUPlugin_dcache_data_load = memaccess_LSUPlugin_dcache_lw;
    end else if((memaccess_MEM_CTRL == MemCtrlEnum_LWU)) begin
        memaccess_LSUPlugin_dcache_data_load = memaccess_LSUPlugin_dcache_lwu;
    end else if((memaccess_MEM_CTRL == MemCtrlEnum_LD)) begin
        memaccess_LSUPlugin_dcache_data_load = memaccess_LSUPlugin_dcache_rdata;
    end else begin
        memaccess_LSUPlugin_dcache_data_load = 64'h0;
    end
  end

  always @(*) begin
    if((memaccess_MEM_CTRL == MemCtrlEnum_LB)) begin
        memaccess_LSUPlugin_lsu_size = 3'b000;
    end else if((memaccess_MEM_CTRL == MemCtrlEnum_LBU)) begin
        memaccess_LSUPlugin_lsu_size = 3'b000;
    end else if((memaccess_MEM_CTRL == MemCtrlEnum_LH)) begin
        memaccess_LSUPlugin_lsu_size = 3'b001;
    end else if((memaccess_MEM_CTRL == MemCtrlEnum_LHU)) begin
        memaccess_LSUPlugin_lsu_size = 3'b001;
    end else if((memaccess_MEM_CTRL == MemCtrlEnum_LW)) begin
        memaccess_LSUPlugin_lsu_size = 3'b010;
    end else if((memaccess_MEM_CTRL == MemCtrlEnum_LWU)) begin
        memaccess_LSUPlugin_lsu_size = 3'b010;
    end else if((memaccess_MEM_CTRL == MemCtrlEnum_LD)) begin
        memaccess_LSUPlugin_lsu_size = 3'b011;
    end else begin
        memaccess_LSUPlugin_lsu_size = 3'b000;
    end
  end

  always @(*) begin
    if((memaccess_MEM_CTRL == MemCtrlEnum_SB)) begin
        memaccess_LSUPlugin_dcache_wdata = memaccess_LSUPlugin_dcache_sb;
    end else if((memaccess_MEM_CTRL == MemCtrlEnum_SH)) begin
        memaccess_LSUPlugin_dcache_wdata = memaccess_LSUPlugin_dcache_sh;
    end else if((memaccess_MEM_CTRL == MemCtrlEnum_SW)) begin
        memaccess_LSUPlugin_dcache_wdata = memaccess_LSUPlugin_dcache_sw;
    end else if((memaccess_MEM_CTRL == MemCtrlEnum_SD)) begin
        memaccess_LSUPlugin_dcache_wdata = memaccess_MEM_WDATA;
    end else begin
        memaccess_LSUPlugin_dcache_wdata = 64'h0;
    end
  end

  assign _zz_4 = zz__zz_memaccess_LSUPlugin_dcache_wstrb(1'b0);
  always @(*) _zz_memaccess_LSUPlugin_dcache_wstrb = _zz_4;
  always @(*) begin
    if((memaccess_MEM_CTRL == MemCtrlEnum_SB)) begin
        memaccess_LSUPlugin_dcache_wstrb = _zz_memaccess_LSUPlugin_dcache_wstrb;
    end else if((memaccess_MEM_CTRL == MemCtrlEnum_SH)) begin
        memaccess_LSUPlugin_dcache_wstrb = _zz_memaccess_LSUPlugin_dcache_wstrb_1;
    end else if((memaccess_MEM_CTRL == MemCtrlEnum_SW)) begin
        memaccess_LSUPlugin_dcache_wstrb = _zz_memaccess_LSUPlugin_dcache_wstrb_2;
    end else if((memaccess_MEM_CTRL == MemCtrlEnum_SD)) begin
        memaccess_LSUPlugin_dcache_wstrb = _zz_memaccess_LSUPlugin_dcache_wstrb_3;
    end else begin
        memaccess_LSUPlugin_dcache_wstrb = 8'h0;
    end
  end

  assign _zz_5 = zz__zz_memaccess_LSUPlugin_dcache_wstrb_1(1'b0);
  always @(*) _zz_memaccess_LSUPlugin_dcache_wstrb_1 = _zz_5;
  assign _zz_6 = zz__zz_memaccess_LSUPlugin_dcache_wstrb_2(1'b0);
  always @(*) _zz_memaccess_LSUPlugin_dcache_wstrb_2 = _zz_6;
  assign _zz_memaccess_LSUPlugin_dcache_wstrb_3[7 : 0] = 8'hff;
  assign memaccess_LSUPlugin_lsu_rdata = memaccess_LSUPlugin_dcache_data_load;
  assign memaccess_LSUPlugin_lsu_wdata = (memaccess_LSUPlugin_dcache_wdata <<< _zz_memaccess_LSUPlugin_lsu_wdata);
  assign memaccess_LSUPlugin_lsu_addr = memaccess_LSUPlugin_cpu_addr;
  assign memaccess_LSUPlugin_lsu_wen = memaccess_IS_STORE;
  assign memaccess_LSUPlugin_lsu_wstrb = (memaccess_LSUPlugin_dcache_wstrb <<< memaccess_LSUPlugin_cpu_addr_offset);
  assign DCachePlugin_dcache_access_cmd_valid = (((! memaccess_LSUPlugin_is_timer) && memaccess_LSUPlugin_is_mem) && memaccess_arbitration_isValid);
  assign DCachePlugin_dcache_access_cmd_payload_addr = memaccess_LSUPlugin_lsu_addr;
  assign DCachePlugin_dcache_access_cmd_payload_wen = memaccess_LSUPlugin_lsu_wen;
  assign DCachePlugin_dcache_access_cmd_payload_wdata = memaccess_LSUPlugin_lsu_wdata;
  assign DCachePlugin_dcache_access_cmd_payload_wstrb = memaccess_LSUPlugin_lsu_wstrb;
  assign DCachePlugin_dcache_access_cmd_payload_size = memaccess_LSUPlugin_lsu_size;
  assign ICachePlugin_icache_access_cmd_ready = iCache_1_cpu_cmd_ready;
  assign ICachePlugin_icache_access_rsp_valid = iCache_1_cpu_rsp_valid;
  assign ICachePlugin_icache_access_rsp_payload_data = iCache_1_cpu_rsp_payload_data;
  assign icache_ar_fire = (icache_ar_valid && icache_ar_ready);
  assign when_ICachePlugin_l141 = (icache_ar_fire && (4'b0000 < ar_len_cnt));
  assign when_ICachePlugin_l149 = (4'b0000 < ar_len_cnt);
  assign icache_ar_fire_1 = (icache_ar_valid && icache_ar_ready);
  assign icache_ar_fire_2 = (icache_ar_valid && icache_ar_ready);
  assign icache_r_ready = 1'b1;
  assign iCache_1_next_level_rsp_valid = (icache_r_valid && (icache_r_payload_id == 2'b00));
  assign DCachePlugin_dcache_access_cmd_ready = dCache_1_cpu_cmd_ready;
  assign DCachePlugin_dcache_access_rsp_valid = dCache_1_cpu_rsp_valid;
  assign DCachePlugin_dcache_access_rsp_payload_data = dCache_1_cpu_rsp_payload_data;
  assign DCachePlugin_dcache_access_stall = dCache_1_stall;
  assign when_DCachePlugin_l265 = (dCache_1_next_level_cmd_valid && (! dCache_1_next_level_cmd_payload_wen));
  assign when_DCachePlugin_l313 = (dCache_1_next_level_cmd_valid && dCache_1_next_level_cmd_payload_wen);
  assign when_DCachePlugin_l267 = (dCache_1_cpu_bypass_cmd_valid && (! dCache_1_cpu_bypass_cmd_payload_wen));
  assign when_DCachePlugin_l233 = (dCache_1_cpu_bypass_cmd_valid && dCache_1_cpu_bypass_cmd_payload_wen);
  assign when_DCachePlugin_l239 = (when_DCachePlugin_l267 || when_DCachePlugin_l233);
  assign when_DCachePlugin_l254 = (when_DCachePlugin_l265 || when_DCachePlugin_l267);
  assign when_DCachePlugin_l258 = (4'b0000 < _zz_when_DCachePlugin_l258);
  assign dcache_ar_fire = (dcache_ar_valid && dcache_ar_ready);
  assign dcache_ar_fire_1 = (dcache_ar_valid && dcache_ar_ready);
  assign when_DCachePlugin_l269 = (dcache_ar_fire_1 && (4'b0000 < _zz_when_DCachePlugin_l258));
  assign dcache_ar_fire_2 = (dcache_ar_valid && dcache_ar_ready);
  assign dcache_r_ready = 1'b1;
  assign when_DCachePlugin_l303 = (when_DCachePlugin_l313 || when_DCachePlugin_l233);
  assign dcache_aw_fire = (dcache_aw_valid && dcache_aw_ready);
  assign when_DCachePlugin_l335 = (when_DCachePlugin_l313 || when_DCachePlugin_l233);
  assign dcache_w_fire = (dcache_w_valid && dcache_w_ready);
  assign dcache_b_ready = 1'b1;
  assign when_DCachePlugin_l349 = (_zz_when_DCachePlugin_l349 == 1'b0);
  assign dcache_aw_fire_1 = (dcache_aw_valid && dcache_aw_ready);
  assign dcache_w_fire_1 = (dcache_w_valid && dcache_w_ready);
  assign when_DCachePlugin_l350 = (dcache_aw_fire_1 && dcache_w_fire_1);
  assign dcache_aw_fire_2 = (dcache_aw_valid && dcache_aw_ready);
  assign dcache_w_fire_2 = (dcache_w_valid && dcache_w_ready);
  assign when_DCachePlugin_l352 = (dcache_aw_fire_2 || dcache_w_fire_2);
  assign dcache_aw_fire_3 = (dcache_aw_valid && dcache_aw_ready);
  assign dcache_w_fire_3 = (dcache_w_valid && dcache_w_ready);
  assign when_DCachePlugin_l357 = (dcache_aw_fire_3 || dcache_w_fire_3);
  assign when_DCachePlugin_l356 = (_zz_when_DCachePlugin_l349 == 1'b1);
  assign dcache_aw_fire_4 = (dcache_aw_valid && dcache_aw_ready);
  assign dcache_w_fire_4 = (dcache_w_valid && dcache_w_ready);
  assign dcache_aw_fire_5 = (dcache_aw_valid && dcache_aw_ready);
  assign dcache_w_fire_5 = (dcache_w_valid && dcache_w_ready);
  assign dCache_1_next_level_rsp_valid = (dCache_1_next_level_cmd_payload_wen ? dcache_b_valid : (dcache_r_valid && (dcache_r_payload_id == 2'b01)));
  assign dCache_1_next_level_rsp_payload_rvalid = (dcache_r_valid && (dcache_r_payload_id == 2'b01));
  assign dCache_1_cpu_bypass_rsp_valid = (_zz_cpu_bypass_rsp_valid_1 ? (_zz_cpu_bypass_rsp_valid ? dcache_b_valid : (dcache_r_valid && (dcache_r_payload_id == 2'b01))) : 1'b0);
  assign when_Pipeline_l127 = (! decode_arbitration_isStuck);
  assign when_Pipeline_l127_1 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_2 = (! memaccess_arbitration_isStuck);
  assign when_Pipeline_l127_3 = (! writeback_arbitration_isStuck);
  assign when_Pipeline_l127_4 = (! decode_arbitration_isStuck);
  assign when_Pipeline_l127_5 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_6 = (! decode_arbitration_isStuck);
  assign when_Pipeline_l127_7 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_8 = (! memaccess_arbitration_isStuck);
  assign when_Pipeline_l127_9 = (! writeback_arbitration_isStuck);
  assign when_Pipeline_l127_10 = (! decode_arbitration_isStuck);
  assign when_Pipeline_l127_11 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_12 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_13 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_14 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_15 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_16 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_17 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_18 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_19 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_20 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_21 = (! memaccess_arbitration_isStuck);
  assign when_Pipeline_l127_22 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_23 = (! memaccess_arbitration_isStuck);
  assign when_Pipeline_l127_24 = (! writeback_arbitration_isStuck);
  assign when_Pipeline_l127_25 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_26 = (! memaccess_arbitration_isStuck);
  assign when_Pipeline_l127_27 = (! writeback_arbitration_isStuck);
  assign when_Pipeline_l127_28 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_29 = (! memaccess_arbitration_isStuck);
  assign when_Pipeline_l127_30 = (! writeback_arbitration_isStuck);
  assign when_Pipeline_l127_31 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_32 = (! memaccess_arbitration_isStuck);
  assign when_Pipeline_l127_33 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_34 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_35 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_36 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_37 = (! memaccess_arbitration_isStuck);
  assign when_Pipeline_l127_38 = (! writeback_arbitration_isStuck);
  assign when_Pipeline_l127_39 = (! memaccess_arbitration_isStuck);
  assign when_Pipeline_l127_40 = (! writeback_arbitration_isStuck);
  assign fetch_arbitration_isFlushed = (({writeback_arbitration_flushNext,{memaccess_arbitration_flushNext,{execute_arbitration_flushNext,decode_arbitration_flushNext}}} != 4'b0000) || ({writeback_arbitration_flushIt,{memaccess_arbitration_flushIt,{execute_arbitration_flushIt,{decode_arbitration_flushIt,fetch_arbitration_flushIt}}}} != 5'h0));
  assign decode_arbitration_isFlushed = (({writeback_arbitration_flushNext,{memaccess_arbitration_flushNext,execute_arbitration_flushNext}} != 3'b000) || ({writeback_arbitration_flushIt,{memaccess_arbitration_flushIt,{execute_arbitration_flushIt,decode_arbitration_flushIt}}} != 4'b0000));
  assign execute_arbitration_isFlushed = (({writeback_arbitration_flushNext,memaccess_arbitration_flushNext} != 2'b00) || ({writeback_arbitration_flushIt,{memaccess_arbitration_flushIt,execute_arbitration_flushIt}} != 3'b000));
  assign memaccess_arbitration_isFlushed = ((writeback_arbitration_flushNext != 1'b0) || ({writeback_arbitration_flushIt,memaccess_arbitration_flushIt} != 2'b00));
  assign writeback_arbitration_isFlushed = (1'b0 || (writeback_arbitration_flushIt != 1'b0));
  assign fetch_arbitration_isStuckByOthers = (fetch_arbitration_haltByOther || ((((1'b0 || decode_arbitration_isStuck) || execute_arbitration_isStuck) || memaccess_arbitration_isStuck) || writeback_arbitration_isStuck));
  assign fetch_arbitration_isStuck = (fetch_arbitration_haltItself || fetch_arbitration_isStuckByOthers);
  assign fetch_arbitration_isMoving = ((! fetch_arbitration_isStuck) && (! fetch_arbitration_removeIt));
  assign fetch_arbitration_isFiring = ((fetch_arbitration_isValid && (! fetch_arbitration_isStuck)) && (! fetch_arbitration_removeIt));
  assign decode_arbitration_isStuckByOthers = (decode_arbitration_haltByOther || (((1'b0 || execute_arbitration_isStuck) || memaccess_arbitration_isStuck) || writeback_arbitration_isStuck));
  assign decode_arbitration_isStuck = (decode_arbitration_haltItself || decode_arbitration_isStuckByOthers);
  assign decode_arbitration_isMoving = ((! decode_arbitration_isStuck) && (! decode_arbitration_removeIt));
  assign decode_arbitration_isFiring = ((decode_arbitration_isValid && (! decode_arbitration_isStuck)) && (! decode_arbitration_removeIt));
  assign execute_arbitration_isStuckByOthers = (execute_arbitration_haltByOther || ((1'b0 || memaccess_arbitration_isStuck) || writeback_arbitration_isStuck));
  assign execute_arbitration_isStuck = (execute_arbitration_haltItself || execute_arbitration_isStuckByOthers);
  assign execute_arbitration_isMoving = ((! execute_arbitration_isStuck) && (! execute_arbitration_removeIt));
  assign execute_arbitration_isFiring = ((execute_arbitration_isValid && (! execute_arbitration_isStuck)) && (! execute_arbitration_removeIt));
  assign memaccess_arbitration_isStuckByOthers = (memaccess_arbitration_haltByOther || (1'b0 || writeback_arbitration_isStuck));
  assign memaccess_arbitration_isStuck = (memaccess_arbitration_haltItself || memaccess_arbitration_isStuckByOthers);
  assign memaccess_arbitration_isMoving = ((! memaccess_arbitration_isStuck) && (! memaccess_arbitration_removeIt));
  assign memaccess_arbitration_isFiring = ((memaccess_arbitration_isValid && (! memaccess_arbitration_isStuck)) && (! memaccess_arbitration_removeIt));
  assign writeback_arbitration_isStuckByOthers = (writeback_arbitration_haltByOther || 1'b0);
  assign writeback_arbitration_isStuck = (writeback_arbitration_haltItself || writeback_arbitration_isStuckByOthers);
  assign writeback_arbitration_isMoving = ((! writeback_arbitration_isStuck) && (! writeback_arbitration_removeIt));
  assign writeback_arbitration_isFiring = ((writeback_arbitration_isValid && (! writeback_arbitration_isStuck)) && (! writeback_arbitration_removeIt));
  assign when_Pipeline_l163 = ((! fetch_arbitration_isStuck) && (! fetch_arbitration_removeIt));
  assign when_Pipeline_l166 = ((! decode_arbitration_isStuck) || decode_arbitration_removeIt);
  assign when_Pipeline_l163_1 = ((! decode_arbitration_isStuck) && (! decode_arbitration_removeIt));
  assign when_Pipeline_l166_1 = ((! execute_arbitration_isStuck) || execute_arbitration_removeIt);
  assign when_Pipeline_l163_2 = ((! execute_arbitration_isStuck) && (! execute_arbitration_removeIt));
  assign when_Pipeline_l166_2 = ((! memaccess_arbitration_isStuck) || memaccess_arbitration_removeIt);
  assign when_Pipeline_l163_3 = ((! memaccess_arbitration_isStuck) && (! memaccess_arbitration_removeIt));
  assign when_Pipeline_l166_3 = ((! writeback_arbitration_isStuck) || writeback_arbitration_removeIt);
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      pc_next <= 64'h0000000030000000;
      fetch_valid <= 1'b0;
      rsp_flush <= 1'b0;
      fetch_state <= IDLE;
      execute_ALUPlugin_branch_history <= 5'h0;
      icache_ar_valid <= 1'b0;
      icache_ar_payload_id <= 2'b00;
      icache_ar_payload_len <= 8'h0;
      icache_ar_payload_size <= 3'b000;
      icache_ar_payload_burst <= 2'b00;
      icache_ar_payload_addr <= 64'h0;
      ar_len_cnt <= 4'b0000;
      _zz_when_DCachePlugin_l349 <= 1'b0;
      _zz_when_DCachePlugin_l258 <= 4'b0000;
      _zz_cpu_bypass_rsp_valid <= 1'b0;
      _zz_cpu_bypass_rsp_valid_1 <= 1'b0;
      dcache_ar_valid <= 1'b0;
      dcache_ar_payload_id <= 2'b00;
      dcache_ar_payload_len <= 8'h0;
      dcache_ar_payload_size <= 3'b000;
      dcache_ar_payload_burst <= 2'b00;
      dcache_ar_payload_addr <= 64'h0;
      dcache_aw_valid <= 1'b0;
      dcache_aw_payload_id <= 2'b00;
      dcache_aw_payload_len <= 8'h0;
      dcache_aw_payload_size <= 3'b000;
      dcache_aw_payload_burst <= 2'b00;
      dcache_aw_payload_addr <= 64'h0;
      dcache_w_valid <= 1'b0;
      dcache_w_payload_data <= 64'h0;
      dcache_w_payload_strb <= 8'h0;
      dcache_w_payload_last <= 1'b0;
      decode_arbitration_isValid <= 1'b0;
      execute_arbitration_isValid <= 1'b0;
      memaccess_arbitration_isValid <= 1'b0;
      writeback_arbitration_isValid <= 1'b0;
    end else begin
      fetch_state <= fetch_state_next;
      if(when_FetchPlugin_l93) begin
        if(when_FetchPlugin_l94) begin
          rsp_flush <= 1'b1;
        end else begin
          if(when_FetchPlugin_l97) begin
            rsp_flush <= 1'b1;
          end else begin
            if(fetch_FetchPlugin_bpu_predict_taken) begin
              rsp_flush <= 1'b1;
            end
          end
        end
      end else begin
        if(ICachePlugin_icache_access_rsp_valid) begin
          rsp_flush <= 1'b0;
        end
      end
      if(when_FetchPlugin_l109) begin
        fetch_valid <= 1'b1;
      end else begin
        fetch_valid <= 1'b0;
      end
      if(when_FetchPlugin_l94) begin
        pc_next <= fetch_INT_PC;
      end else begin
        if(when_FetchPlugin_l97) begin
          pc_next <= _zz_pc_next;
        end else begin
          if(fetch_FetchPlugin_bpu_predict_taken) begin
            pc_next <= fetch_BPU_PC_NEXT;
          end else begin
            if(ICachePlugin_icache_access_cmd_fire_1) begin
              pc_next <= (pc_next + 64'h0000000000000004);
            end
          end
        end
      end
      if(execute_arbitration_isFiring) begin
        execute_ALUPlugin_branch_history <= {execute_ALUPlugin_branch_history[3 : 0],execute_ALUPlugin_branch_taken};
      end
      if(iCache_1_next_level_cmd_valid) begin
        ar_len_cnt <= iCache_1_next_level_cmd_payload_len;
      end else begin
        if(when_ICachePlugin_l141) begin
          ar_len_cnt <= (ar_len_cnt - 4'b0001);
        end
      end
      if(iCache_1_next_level_cmd_valid) begin
        icache_ar_valid <= 1'b1;
      end else begin
        if(icache_ar_fire_1) begin
          if(when_ICachePlugin_l149) begin
            icache_ar_valid <= 1'b1;
          end else begin
            icache_ar_valid <= 1'b0;
          end
        end
      end
      icache_ar_payload_id <= 2'b00;
      icache_ar_payload_len <= 8'h0;
      icache_ar_payload_size <= iCache_1_next_level_cmd_payload_size;
      icache_ar_payload_burst <= 2'b01;
      if(iCache_1_next_level_cmd_valid) begin
        icache_ar_payload_addr <= iCache_1_next_level_cmd_payload_addr;
      end else begin
        if(icache_ar_fire_2) begin
          icache_ar_payload_addr <= (icache_ar_payload_addr + 64'h0000000000000008);
        end
      end
      if(when_DCachePlugin_l233) begin
        _zz_cpu_bypass_rsp_valid <= 1'b1;
      end else begin
        if(dCache_1_cpu_bypass_rsp_valid) begin
          _zz_cpu_bypass_rsp_valid <= 1'b0;
        end
      end
      if(when_DCachePlugin_l239) begin
        _zz_cpu_bypass_rsp_valid_1 <= 1'b1;
      end else begin
        if(dCache_1_cpu_bypass_rsp_valid) begin
          _zz_cpu_bypass_rsp_valid_1 <= 1'b0;
        end
      end
      if(when_DCachePlugin_l254) begin
        dcache_ar_valid <= 1'b1;
      end else begin
        if(dcache_ar_fire) begin
          if(when_DCachePlugin_l258) begin
            dcache_ar_valid <= 1'b1;
          end else begin
            dcache_ar_valid <= 1'b0;
          end
        end
      end
      if(when_DCachePlugin_l265) begin
        _zz_when_DCachePlugin_l258 <= dCache_1_next_level_cmd_payload_len;
      end else begin
        if(when_DCachePlugin_l267) begin
          _zz_when_DCachePlugin_l258 <= 4'b0000;
        end else begin
          if(when_DCachePlugin_l269) begin
            _zz_when_DCachePlugin_l258 <= (_zz_when_DCachePlugin_l258 - 4'b0001);
          end
        end
      end
      dcache_ar_payload_id <= 2'b01;
      dcache_ar_payload_len <= 8'h0;
      if(when_DCachePlugin_l267) begin
        dcache_ar_payload_size <= dCache_1_cpu_bypass_cmd_payload_size;
      end else begin
        if(dCache_1_next_level_cmd_valid) begin
          dcache_ar_payload_size <= dCache_1_next_level_cmd_payload_size;
        end
      end
      dcache_ar_payload_burst <= 2'b01;
      if(when_DCachePlugin_l265) begin
        dcache_ar_payload_addr <= dCache_1_next_level_cmd_payload_addr;
      end else begin
        if(when_DCachePlugin_l267) begin
          dcache_ar_payload_addr <= dCache_1_cpu_bypass_cmd_payload_addr;
        end else begin
          if(dcache_ar_fire_2) begin
            dcache_ar_payload_addr <= (dcache_ar_payload_addr + 64'h0000000000000008);
          end
        end
      end
      if(when_DCachePlugin_l303) begin
        dcache_aw_valid <= 1'b1;
      end else begin
        if(dcache_aw_fire) begin
          dcache_aw_valid <= 1'b0;
        end
      end
      dcache_aw_payload_id <= 2'b10;
      if(when_DCachePlugin_l233) begin
        dcache_aw_payload_len <= 8'h0;
      end else begin
        if(when_DCachePlugin_l313) begin
          dcache_aw_payload_len <= {4'd0, dCache_1_next_level_cmd_payload_len};
        end
      end
      if(when_DCachePlugin_l233) begin
        dcache_aw_payload_size <= dCache_1_cpu_bypass_cmd_payload_size;
      end else begin
        if(when_DCachePlugin_l313) begin
          dcache_aw_payload_size <= dCache_1_next_level_cmd_payload_size;
        end
      end
      dcache_aw_payload_burst <= 2'b01;
      if(when_DCachePlugin_l233) begin
        dcache_aw_payload_addr <= dCache_1_cpu_bypass_cmd_payload_addr;
      end else begin
        if(when_DCachePlugin_l313) begin
          dcache_aw_payload_addr <= dCache_1_next_level_cmd_payload_addr;
        end
      end
      if(when_DCachePlugin_l335) begin
        dcache_w_valid <= 1'b1;
      end else begin
        if(dcache_w_fire) begin
          dcache_w_valid <= 1'b0;
        end
      end
      dcache_w_payload_data <= (when_DCachePlugin_l233 ? dCache_1_cpu_bypass_cmd_payload_wdata : dCache_1_next_level_cmd_payload_wdata);
      dcache_w_payload_strb <= (when_DCachePlugin_l233 ? dCache_1_cpu_bypass_cmd_payload_wstrb : dCache_1_next_level_cmd_payload_wstrb);
      dcache_w_payload_last <= 1'b1;
      if(when_DCachePlugin_l349) begin
        if(when_DCachePlugin_l350) begin
          _zz_when_DCachePlugin_l349 <= 1'b0;
        end else begin
          if(when_DCachePlugin_l352) begin
            _zz_when_DCachePlugin_l349 <= 1'b1;
          end
        end
      end else begin
        if(when_DCachePlugin_l356) begin
          if(when_DCachePlugin_l357) begin
            _zz_when_DCachePlugin_l349 <= 1'b0;
          end
        end
      end
      if(when_Pipeline_l163) begin
        decode_arbitration_isValid <= fetch_arbitration_isValid;
      end else begin
        if(when_Pipeline_l166) begin
          decode_arbitration_isValid <= 1'b0;
        end
      end
      if(when_Pipeline_l163_1) begin
        execute_arbitration_isValid <= decode_arbitration_isValid;
      end else begin
        if(when_Pipeline_l166_1) begin
          execute_arbitration_isValid <= 1'b0;
        end
      end
      if(when_Pipeline_l163_2) begin
        memaccess_arbitration_isValid <= execute_arbitration_isValid;
      end else begin
        if(when_Pipeline_l166_2) begin
          memaccess_arbitration_isValid <= 1'b0;
        end
      end
      if(when_Pipeline_l163_3) begin
        writeback_arbitration_isValid <= memaccess_arbitration_isValid;
      end else begin
        if(when_Pipeline_l166_3) begin
          writeback_arbitration_isValid <= 1'b0;
        end
      end
    end
  end

  always @(posedge io_axiClk) begin
    if(when_Pipeline_l127) begin
      fetch_to_decode_PC <= fetch_PC;
    end
    if(when_Pipeline_l127_1) begin
      decode_to_execute_PC <= decode_PC;
    end
    if(when_Pipeline_l127_2) begin
      execute_to_memaccess_PC <= _zz_execute_to_memaccess_PC;
    end
    if(when_Pipeline_l127_3) begin
      memaccess_to_writeback_PC <= memaccess_PC;
    end
    if(when_Pipeline_l127_4) begin
      fetch_to_decode_PC_NEXT <= fetch_PC_NEXT;
    end
    if(when_Pipeline_l127_5) begin
      decode_to_execute_PC_NEXT <= decode_PC_NEXT;
    end
    if(when_Pipeline_l127_6) begin
      fetch_to_decode_INSTRUCTION <= fetch_INSTRUCTION;
    end
    if(when_Pipeline_l127_7) begin
      decode_to_execute_INSTRUCTION <= decode_INSTRUCTION;
    end
    if(when_Pipeline_l127_8) begin
      execute_to_memaccess_INSTRUCTION <= execute_INSTRUCTION;
    end
    if(when_Pipeline_l127_9) begin
      memaccess_to_writeback_INSTRUCTION <= memaccess_INSTRUCTION;
    end
    if(when_Pipeline_l127_10) begin
      fetch_to_decode_PREDICT_TAKEN <= fetch_PREDICT_TAKEN;
    end
    if(when_Pipeline_l127_11) begin
      decode_to_execute_PREDICT_TAKEN <= decode_PREDICT_TAKEN;
    end
    if(when_Pipeline_l127_12) begin
      decode_to_execute_IMM <= decode_IMM;
    end
    if(when_Pipeline_l127_13) begin
      decode_to_execute_RS1 <= decode_RS1;
    end
    if(when_Pipeline_l127_14) begin
      decode_to_execute_RS2 <= decode_RS2;
    end
    if(when_Pipeline_l127_15) begin
      decode_to_execute_RS1_ADDR <= decode_RS1_ADDR;
    end
    if(when_Pipeline_l127_16) begin
      decode_to_execute_RS2_ADDR <= decode_RS2_ADDR;
    end
    if(when_Pipeline_l127_17) begin
      decode_to_execute_ALU_CTRL <= decode_ALU_CTRL;
    end
    if(when_Pipeline_l127_18) begin
      decode_to_execute_ALU_WORD <= decode_ALU_WORD;
    end
    if(when_Pipeline_l127_19) begin
      decode_to_execute_SRC2_IS_IMM <= decode_SRC2_IS_IMM;
    end
    if(when_Pipeline_l127_20) begin
      decode_to_execute_MEM_CTRL <= decode_MEM_CTRL;
    end
    if(when_Pipeline_l127_21) begin
      execute_to_memaccess_MEM_CTRL <= execute_MEM_CTRL;
    end
    if(when_Pipeline_l127_22) begin
      decode_to_execute_RD_WEN <= decode_RD_WEN;
    end
    if(when_Pipeline_l127_23) begin
      execute_to_memaccess_RD_WEN <= execute_RD_WEN;
    end
    if(when_Pipeline_l127_24) begin
      memaccess_to_writeback_RD_WEN <= _zz_DecodePlugin_hazard_rs1_from_mem_3;
    end
    if(when_Pipeline_l127_25) begin
      decode_to_execute_RD_ADDR <= decode_RD_ADDR;
    end
    if(when_Pipeline_l127_26) begin
      execute_to_memaccess_RD_ADDR <= execute_RD_ADDR;
    end
    if(when_Pipeline_l127_27) begin
      memaccess_to_writeback_RD_ADDR <= _zz_DecodePlugin_hazard_rs1_from_mem_2;
    end
    if(when_Pipeline_l127_28) begin
      decode_to_execute_IS_LOAD <= decode_IS_LOAD;
    end
    if(when_Pipeline_l127_29) begin
      execute_to_memaccess_IS_LOAD <= execute_IS_LOAD;
    end
    if(when_Pipeline_l127_30) begin
      memaccess_to_writeback_IS_LOAD <= _zz_DecodePlugin_hazard_rs1_from_mem;
    end
    if(when_Pipeline_l127_31) begin
      decode_to_execute_IS_STORE <= decode_IS_STORE;
    end
    if(when_Pipeline_l127_32) begin
      execute_to_memaccess_IS_STORE <= execute_IS_STORE;
    end
    if(when_Pipeline_l127_33) begin
      decode_to_execute_CSR_CTRL <= decode_CSR_CTRL;
    end
    if(when_Pipeline_l127_34) begin
      decode_to_execute_CSR_ADDR <= _zz_decode_to_execute_CSR_ADDR;
    end
    if(when_Pipeline_l127_35) begin
      decode_to_execute_CSR_WEN <= decode_CSR_WEN;
    end
    if(when_Pipeline_l127_36) begin
      decode_to_execute_CSR_RDATA <= decode_CSR_RDATA;
    end
    if(when_Pipeline_l127_37) begin
      execute_to_memaccess_ALU_RESULT <= execute_ALU_RESULT;
    end
    if(when_Pipeline_l127_38) begin
      memaccess_to_writeback_ALU_RESULT <= _zz_execute_MEM_WDATA_1;
    end
    if(when_Pipeline_l127_39) begin
      execute_to_memaccess_MEM_WDATA <= execute_MEM_WDATA;
    end
    if(when_Pipeline_l127_40) begin
      memaccess_to_writeback_LSU_RDATA <= _zz_execute_MEM_WDATA;
    end
  end


endmodule

module BufferCC (
  input               io_dataIn,
  output              io_dataOut,
  input               io_axiClk,
  input               io_asyncResetn
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_axiClk) begin
    buffers_0 <= io_dataIn;
    buffers_1 <= buffers_0;
  end


endmodule

//StreamFifoLowLatency replaced by StreamFifoLowLatency_2

module StreamArbiter (
  input               io_inputs_0_valid,
  output              io_inputs_0_ready,
  input      [19:0]   io_inputs_0_payload_addr,
  input      [3:0]    io_inputs_0_payload_id,
  input      [7:0]    io_inputs_0_payload_len,
  input      [2:0]    io_inputs_0_payload_size,
  input      [1:0]    io_inputs_0_payload_burst,
  input               io_inputs_0_payload_write,
  input               io_inputs_1_valid,
  output              io_inputs_1_ready,
  input      [19:0]   io_inputs_1_payload_addr,
  input      [3:0]    io_inputs_1_payload_id,
  input      [7:0]    io_inputs_1_payload_len,
  input      [2:0]    io_inputs_1_payload_size,
  input      [1:0]    io_inputs_1_payload_burst,
  input               io_inputs_1_payload_write,
  output              io_output_valid,
  input               io_output_ready,
  output     [19:0]   io_output_payload_addr,
  output     [3:0]    io_output_payload_id,
  output     [7:0]    io_output_payload_len,
  output     [2:0]    io_output_payload_size,
  output     [1:0]    io_output_payload_burst,
  output              io_output_payload_write,
  output     [0:0]    io_chosen,
  output     [1:0]    io_chosenOH,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  wire       [3:0]    _zz__zz_maskProposal_0_2;
  wire       [3:0]    _zz__zz_maskProposal_0_2_1;
  wire       [1:0]    _zz__zz_maskProposal_0_2_2;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire       [1:0]    _zz_maskProposal_0;
  wire       [3:0]    _zz_maskProposal_0_1;
  wire       [3:0]    _zz_maskProposal_0_2;
  wire       [1:0]    _zz_maskProposal_0_3;
  wire                io_output_fire;
  wire                _zz_io_chosen;

  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = {maskLocked_0,maskLocked_1};
  assign _zz__zz_maskProposal_0_2_1 = {2'd0, _zz__zz_maskProposal_0_2_2};
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign _zz_maskProposal_0 = {io_inputs_1_valid,io_inputs_0_valid};
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[3 : 2] | _zz_maskProposal_0_2[1 : 0]);
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign maskProposal_1 = _zz_maskProposal_0_3[1];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_valid = ((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1));
  assign io_output_payload_addr = (maskRouted_0 ? io_inputs_0_payload_addr : io_inputs_1_payload_addr);
  assign io_output_payload_id = (maskRouted_0 ? io_inputs_0_payload_id : io_inputs_1_payload_id);
  assign io_output_payload_len = (maskRouted_0 ? io_inputs_0_payload_len : io_inputs_1_payload_len);
  assign io_output_payload_size = (maskRouted_0 ? io_inputs_0_payload_size : io_inputs_1_payload_size);
  assign io_output_payload_burst = (maskRouted_0 ? io_inputs_0_payload_burst : io_inputs_1_payload_burst);
  assign io_output_payload_write = (maskRouted_0 ? io_inputs_0_payload_write : io_inputs_1_payload_write);
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_chosenOH = {maskRouted_1,maskRouted_0};
  assign _zz_io_chosen = io_chosenOH[1];
  assign io_chosen = _zz_io_chosen;
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b0;
      maskLocked_1 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

//StreamFifoLowLatency_1 replaced by StreamFifoLowLatency_2

module StreamArbiter_1 (
  input               io_inputs_0_valid,
  output              io_inputs_0_ready,
  input      [16:0]   io_inputs_0_payload_addr,
  input      [3:0]    io_inputs_0_payload_id,
  input      [7:0]    io_inputs_0_payload_len,
  input      [2:0]    io_inputs_0_payload_size,
  input      [1:0]    io_inputs_0_payload_burst,
  input               io_inputs_0_payload_write,
  input               io_inputs_1_valid,
  output              io_inputs_1_ready,
  input      [16:0]   io_inputs_1_payload_addr,
  input      [3:0]    io_inputs_1_payload_id,
  input      [7:0]    io_inputs_1_payload_len,
  input      [2:0]    io_inputs_1_payload_size,
  input      [1:0]    io_inputs_1_payload_burst,
  input               io_inputs_1_payload_write,
  output              io_output_valid,
  input               io_output_ready,
  output     [16:0]   io_output_payload_addr,
  output     [3:0]    io_output_payload_id,
  output     [7:0]    io_output_payload_len,
  output     [2:0]    io_output_payload_size,
  output     [1:0]    io_output_payload_burst,
  output              io_output_payload_write,
  output     [0:0]    io_chosen,
  output     [1:0]    io_chosenOH,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  wire       [3:0]    _zz__zz_maskProposal_0_2;
  wire       [3:0]    _zz__zz_maskProposal_0_2_1;
  wire       [1:0]    _zz__zz_maskProposal_0_2_2;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire       [1:0]    _zz_maskProposal_0;
  wire       [3:0]    _zz_maskProposal_0_1;
  wire       [3:0]    _zz_maskProposal_0_2;
  wire       [1:0]    _zz_maskProposal_0_3;
  wire                io_output_fire;
  wire                _zz_io_chosen;

  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = {maskLocked_0,maskLocked_1};
  assign _zz__zz_maskProposal_0_2_1 = {2'd0, _zz__zz_maskProposal_0_2_2};
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign _zz_maskProposal_0 = {io_inputs_1_valid,io_inputs_0_valid};
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[3 : 2] | _zz_maskProposal_0_2[1 : 0]);
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign maskProposal_1 = _zz_maskProposal_0_3[1];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_valid = ((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1));
  assign io_output_payload_addr = (maskRouted_0 ? io_inputs_0_payload_addr : io_inputs_1_payload_addr);
  assign io_output_payload_id = (maskRouted_0 ? io_inputs_0_payload_id : io_inputs_1_payload_id);
  assign io_output_payload_len = (maskRouted_0 ? io_inputs_0_payload_len : io_inputs_1_payload_len);
  assign io_output_payload_size = (maskRouted_0 ? io_inputs_0_payload_size : io_inputs_1_payload_size);
  assign io_output_payload_burst = (maskRouted_0 ? io_inputs_0_payload_burst : io_inputs_1_payload_burst);
  assign io_output_payload_write = (maskRouted_0 ? io_inputs_0_payload_write : io_inputs_1_payload_write);
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_chosenOH = {maskRouted_1,maskRouted_0};
  assign _zz_io_chosen = io_chosenOH[1];
  assign io_chosen = _zz_io_chosen;
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b0;
      maskLocked_1 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

module Axi4WriteOnlyErrorSlave (
  input               io_axi_aw_valid,
  output              io_axi_aw_ready,
  input      [31:0]   io_axi_aw_payload_addr,
  input      [3:0]    io_axi_aw_payload_id,
  input      [3:0]    io_axi_aw_payload_region,
  input      [7:0]    io_axi_aw_payload_len,
  input      [2:0]    io_axi_aw_payload_size,
  input      [1:0]    io_axi_aw_payload_burst,
  input      [0:0]    io_axi_aw_payload_lock,
  input      [3:0]    io_axi_aw_payload_cache,
  input      [3:0]    io_axi_aw_payload_qos,
  input      [2:0]    io_axi_aw_payload_prot,
  input               io_axi_w_valid,
  output              io_axi_w_ready,
  input      [31:0]   io_axi_w_payload_data,
  input      [3:0]    io_axi_w_payload_strb,
  input               io_axi_w_payload_last,
  output              io_axi_b_valid,
  input               io_axi_b_ready,
  output     [3:0]    io_axi_b_payload_id,
  output     [1:0]    io_axi_b_payload_resp,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  reg                 consumeData;
  reg                 sendRsp;
  reg        [3:0]    id;
  wire                io_axi_aw_fire;
  wire                io_axi_w_fire;
  wire                when_Axi4ErrorSlave_l24;
  wire                io_axi_b_fire;

  assign io_axi_aw_ready = (! (consumeData || sendRsp));
  assign io_axi_aw_fire = (io_axi_aw_valid && io_axi_aw_ready);
  assign io_axi_w_ready = consumeData;
  assign io_axi_w_fire = (io_axi_w_valid && io_axi_w_ready);
  assign when_Axi4ErrorSlave_l24 = (io_axi_w_fire && io_axi_w_payload_last);
  assign io_axi_b_valid = sendRsp;
  assign io_axi_b_payload_resp = 2'b11;
  assign io_axi_b_payload_id = id;
  assign io_axi_b_fire = (io_axi_b_valid && io_axi_b_ready);
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      consumeData <= 1'b0;
      sendRsp <= 1'b0;
    end else begin
      if(io_axi_aw_fire) begin
        consumeData <= 1'b1;
      end
      if(when_Axi4ErrorSlave_l24) begin
        consumeData <= 1'b0;
        sendRsp <= 1'b1;
      end
      if(io_axi_b_fire) begin
        sendRsp <= 1'b0;
      end
    end
  end

  always @(posedge io_axiClk) begin
    if(io_axi_aw_fire) begin
      id <= io_axi_aw_payload_id;
    end
  end


endmodule

module Axi4ReadOnlyErrorSlave (
  input               io_axi_ar_valid,
  output              io_axi_ar_ready,
  input      [31:0]   io_axi_ar_payload_addr,
  input      [3:0]    io_axi_ar_payload_id,
  input      [3:0]    io_axi_ar_payload_region,
  input      [7:0]    io_axi_ar_payload_len,
  input      [2:0]    io_axi_ar_payload_size,
  input      [1:0]    io_axi_ar_payload_burst,
  input      [0:0]    io_axi_ar_payload_lock,
  input      [3:0]    io_axi_ar_payload_cache,
  input      [3:0]    io_axi_ar_payload_qos,
  input      [2:0]    io_axi_ar_payload_prot,
  output              io_axi_r_valid,
  input               io_axi_r_ready,
  output     [31:0]   io_axi_r_payload_data,
  output     [3:0]    io_axi_r_payload_id,
  output     [1:0]    io_axi_r_payload_resp,
  output              io_axi_r_payload_last,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  reg                 sendRsp;
  reg        [3:0]    id;
  reg        [7:0]    remaining;
  wire                remainingZero;
  wire                io_axi_ar_fire;

  assign remainingZero = (remaining == 8'h0);
  assign io_axi_ar_ready = (! sendRsp);
  assign io_axi_ar_fire = (io_axi_ar_valid && io_axi_ar_ready);
  assign io_axi_r_valid = sendRsp;
  assign io_axi_r_payload_id = id;
  assign io_axi_r_payload_resp = 2'b11;
  assign io_axi_r_payload_last = remainingZero;
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      sendRsp <= 1'b0;
    end else begin
      if(io_axi_ar_fire) begin
        sendRsp <= 1'b1;
      end
      if(sendRsp) begin
        if(io_axi_r_ready) begin
          if(remainingZero) begin
            sendRsp <= 1'b0;
          end
        end
      end
    end
  end

  always @(posedge io_axiClk) begin
    if(io_axi_ar_fire) begin
      remaining <= io_axi_ar_payload_len;
      id <= io_axi_ar_payload_id;
    end
    if(sendRsp) begin
      if(io_axi_r_ready) begin
        remaining <= (remaining - 8'h01);
      end
    end
  end


endmodule

module StreamArbiter_2 (
  input               io_inputs_0_valid,
  output              io_inputs_0_ready,
  input      [31:0]   io_inputs_0_payload_addr,
  input      [2:0]    io_inputs_0_payload_id,
  input      [3:0]    io_inputs_0_payload_region,
  input      [7:0]    io_inputs_0_payload_len,
  input      [2:0]    io_inputs_0_payload_size,
  input      [1:0]    io_inputs_0_payload_burst,
  input      [0:0]    io_inputs_0_payload_lock,
  input      [3:0]    io_inputs_0_payload_cache,
  input      [3:0]    io_inputs_0_payload_qos,
  input      [2:0]    io_inputs_0_payload_prot,
  input               io_inputs_1_valid,
  output              io_inputs_1_ready,
  input      [31:0]   io_inputs_1_payload_addr,
  input      [2:0]    io_inputs_1_payload_id,
  input      [3:0]    io_inputs_1_payload_region,
  input      [7:0]    io_inputs_1_payload_len,
  input      [2:0]    io_inputs_1_payload_size,
  input      [1:0]    io_inputs_1_payload_burst,
  input      [0:0]    io_inputs_1_payload_lock,
  input      [3:0]    io_inputs_1_payload_cache,
  input      [3:0]    io_inputs_1_payload_qos,
  input      [2:0]    io_inputs_1_payload_prot,
  output              io_output_valid,
  input               io_output_ready,
  output     [31:0]   io_output_payload_addr,
  output     [2:0]    io_output_payload_id,
  output     [3:0]    io_output_payload_region,
  output     [7:0]    io_output_payload_len,
  output     [2:0]    io_output_payload_size,
  output     [1:0]    io_output_payload_burst,
  output     [0:0]    io_output_payload_lock,
  output     [3:0]    io_output_payload_cache,
  output     [3:0]    io_output_payload_qos,
  output     [2:0]    io_output_payload_prot,
  output     [0:0]    io_chosen,
  output     [1:0]    io_chosenOH,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  wire       [3:0]    _zz__zz_maskProposal_0_2;
  wire       [3:0]    _zz__zz_maskProposal_0_2_1;
  wire       [1:0]    _zz__zz_maskProposal_0_2_2;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire       [1:0]    _zz_maskProposal_0;
  wire       [3:0]    _zz_maskProposal_0_1;
  wire       [3:0]    _zz_maskProposal_0_2;
  wire       [1:0]    _zz_maskProposal_0_3;
  wire                io_output_fire;
  wire                _zz_io_chosen;

  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = {maskLocked_0,maskLocked_1};
  assign _zz__zz_maskProposal_0_2_1 = {2'd0, _zz__zz_maskProposal_0_2_2};
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign _zz_maskProposal_0 = {io_inputs_1_valid,io_inputs_0_valid};
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[3 : 2] | _zz_maskProposal_0_2[1 : 0]);
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign maskProposal_1 = _zz_maskProposal_0_3[1];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_valid = ((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1));
  assign io_output_payload_addr = (maskRouted_0 ? io_inputs_0_payload_addr : io_inputs_1_payload_addr);
  assign io_output_payload_id = (maskRouted_0 ? io_inputs_0_payload_id : io_inputs_1_payload_id);
  assign io_output_payload_region = (maskRouted_0 ? io_inputs_0_payload_region : io_inputs_1_payload_region);
  assign io_output_payload_len = (maskRouted_0 ? io_inputs_0_payload_len : io_inputs_1_payload_len);
  assign io_output_payload_size = (maskRouted_0 ? io_inputs_0_payload_size : io_inputs_1_payload_size);
  assign io_output_payload_burst = (maskRouted_0 ? io_inputs_0_payload_burst : io_inputs_1_payload_burst);
  assign io_output_payload_lock = (maskRouted_0 ? io_inputs_0_payload_lock : io_inputs_1_payload_lock);
  assign io_output_payload_cache = (maskRouted_0 ? io_inputs_0_payload_cache : io_inputs_1_payload_cache);
  assign io_output_payload_qos = (maskRouted_0 ? io_inputs_0_payload_qos : io_inputs_1_payload_qos);
  assign io_output_payload_prot = (maskRouted_0 ? io_inputs_0_payload_prot : io_inputs_1_payload_prot);
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_chosenOH = {maskRouted_1,maskRouted_0};
  assign _zz_io_chosen = io_chosenOH[1];
  assign io_chosen = _zz_io_chosen;
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b0;
      maskLocked_1 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

module StreamFifoLowLatency_2 (
  input               io_push_valid,
  output              io_push_ready,
  output reg          io_pop_valid,
  input               io_pop_ready,
  input               io_flush,
  output     [2:0]    io_occupancy,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  wire       [1:0]    _zz_pushPtr_valueNext;
  wire       [0:0]    _zz_pushPtr_valueNext_1;
  wire       [1:0]    _zz_popPtr_valueNext;
  wire       [0:0]    _zz_popPtr_valueNext_1;
  reg                 pushPtr_willIncrement;
  reg                 pushPtr_willClear;
  reg        [1:0]    pushPtr_valueNext;
  reg        [1:0]    pushPtr_value;
  wire                pushPtr_willOverflowIfInc;
  wire                pushPtr_willOverflow;
  reg                 popPtr_willIncrement;
  reg                 popPtr_willClear;
  reg        [1:0]    popPtr_valueNext;
  reg        [1:0]    popPtr_value;
  wire                popPtr_willOverflowIfInc;
  wire                popPtr_willOverflow;
  wire                ptrMatch;
  reg                 risingOccupancy;
  wire                empty;
  wire                full;
  wire                pushing;
  wire                popping;
  wire                when_Stream_l1217;
  wire                when_Stream_l1230;
  wire       [1:0]    ptrDif;

  assign _zz_pushPtr_valueNext_1 = pushPtr_willIncrement;
  assign _zz_pushPtr_valueNext = {1'd0, _zz_pushPtr_valueNext_1};
  assign _zz_popPtr_valueNext_1 = popPtr_willIncrement;
  assign _zz_popPtr_valueNext = {1'd0, _zz_popPtr_valueNext_1};
  always @(*) begin
    pushPtr_willIncrement = 1'b0;
    if(pushing) begin
      pushPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    pushPtr_willClear = 1'b0;
    if(io_flush) begin
      pushPtr_willClear = 1'b1;
    end
  end

  assign pushPtr_willOverflowIfInc = (pushPtr_value == 2'b11);
  assign pushPtr_willOverflow = (pushPtr_willOverflowIfInc && pushPtr_willIncrement);
  always @(*) begin
    pushPtr_valueNext = (pushPtr_value + _zz_pushPtr_valueNext);
    if(pushPtr_willClear) begin
      pushPtr_valueNext = 2'b00;
    end
  end

  always @(*) begin
    popPtr_willIncrement = 1'b0;
    if(popping) begin
      popPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    popPtr_willClear = 1'b0;
    if(io_flush) begin
      popPtr_willClear = 1'b1;
    end
  end

  assign popPtr_willOverflowIfInc = (popPtr_value == 2'b11);
  assign popPtr_willOverflow = (popPtr_willOverflowIfInc && popPtr_willIncrement);
  always @(*) begin
    popPtr_valueNext = (popPtr_value + _zz_popPtr_valueNext);
    if(popPtr_willClear) begin
      popPtr_valueNext = 2'b00;
    end
  end

  assign ptrMatch = (pushPtr_value == popPtr_value);
  assign empty = (ptrMatch && (! risingOccupancy));
  assign full = (ptrMatch && risingOccupancy);
  assign pushing = (io_push_valid && io_push_ready);
  assign popping = (io_pop_valid && io_pop_ready);
  assign io_push_ready = (! full);
  assign when_Stream_l1217 = (! empty);
  always @(*) begin
    if(when_Stream_l1217) begin
      io_pop_valid = 1'b1;
    end else begin
      io_pop_valid = io_push_valid;
    end
  end

  assign when_Stream_l1230 = (pushing != popping);
  assign ptrDif = (pushPtr_value - popPtr_value);
  assign io_occupancy = {(risingOccupancy && ptrMatch),ptrDif};
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      pushPtr_value <= 2'b00;
      popPtr_value <= 2'b00;
      risingOccupancy <= 1'b0;
    end else begin
      pushPtr_value <= pushPtr_valueNext;
      popPtr_value <= popPtr_valueNext;
      if(when_Stream_l1230) begin
        risingOccupancy <= pushing;
      end
      if(io_flush) begin
        risingOccupancy <= 1'b0;
      end
    end
  end


endmodule

module StreamArbiter_3 (
  input               io_inputs_0_valid,
  output              io_inputs_0_ready,
  input      [16:0]   io_inputs_0_payload_addr,
  input      [2:0]    io_inputs_0_payload_id,
  input      [7:0]    io_inputs_0_payload_len,
  input      [2:0]    io_inputs_0_payload_size,
  input      [1:0]    io_inputs_0_payload_burst,
  input               io_inputs_0_payload_write,
  input               io_inputs_1_valid,
  output              io_inputs_1_ready,
  input      [16:0]   io_inputs_1_payload_addr,
  input      [2:0]    io_inputs_1_payload_id,
  input      [7:0]    io_inputs_1_payload_len,
  input      [2:0]    io_inputs_1_payload_size,
  input      [1:0]    io_inputs_1_payload_burst,
  input               io_inputs_1_payload_write,
  input               io_inputs_2_valid,
  output              io_inputs_2_ready,
  input      [16:0]   io_inputs_2_payload_addr,
  input      [2:0]    io_inputs_2_payload_id,
  input      [7:0]    io_inputs_2_payload_len,
  input      [2:0]    io_inputs_2_payload_size,
  input      [1:0]    io_inputs_2_payload_burst,
  input               io_inputs_2_payload_write,
  output              io_output_valid,
  input               io_output_ready,
  output     [16:0]   io_output_payload_addr,
  output     [2:0]    io_output_payload_id,
  output     [7:0]    io_output_payload_len,
  output     [2:0]    io_output_payload_size,
  output     [1:0]    io_output_payload_burst,
  output              io_output_payload_write,
  output     [1:0]    io_chosen,
  output     [2:0]    io_chosenOH,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  wire       [5:0]    _zz__zz_maskProposal_0_2;
  wire       [5:0]    _zz__zz_maskProposal_0_2_1;
  wire       [2:0]    _zz__zz_maskProposal_0_2_2;
  reg        [16:0]   _zz_io_output_payload_addr_1;
  reg        [2:0]    _zz_io_output_payload_id;
  reg        [7:0]    _zz_io_output_payload_len;
  reg        [2:0]    _zz_io_output_payload_size;
  reg        [1:0]    _zz_io_output_payload_burst;
  reg                 _zz_io_output_payload_write;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  wire                maskProposal_2;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  reg                 maskLocked_2;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire                maskRouted_2;
  wire       [2:0]    _zz_maskProposal_0;
  wire       [5:0]    _zz_maskProposal_0_1;
  wire       [5:0]    _zz_maskProposal_0_2;
  wire       [2:0]    _zz_maskProposal_0_3;
  wire                io_output_fire;
  wire       [1:0]    _zz_io_output_payload_addr;
  wire                _zz_io_chosen;
  wire                _zz_io_chosen_1;

  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = {maskLocked_1,{maskLocked_0,maskLocked_2}};
  assign _zz__zz_maskProposal_0_2_1 = {3'd0, _zz__zz_maskProposal_0_2_2};
  always @(*) begin
    case(_zz_io_output_payload_addr)
      2'b00 : begin
        _zz_io_output_payload_addr_1 = io_inputs_0_payload_addr;
        _zz_io_output_payload_id = io_inputs_0_payload_id;
        _zz_io_output_payload_len = io_inputs_0_payload_len;
        _zz_io_output_payload_size = io_inputs_0_payload_size;
        _zz_io_output_payload_burst = io_inputs_0_payload_burst;
        _zz_io_output_payload_write = io_inputs_0_payload_write;
      end
      2'b01 : begin
        _zz_io_output_payload_addr_1 = io_inputs_1_payload_addr;
        _zz_io_output_payload_id = io_inputs_1_payload_id;
        _zz_io_output_payload_len = io_inputs_1_payload_len;
        _zz_io_output_payload_size = io_inputs_1_payload_size;
        _zz_io_output_payload_burst = io_inputs_1_payload_burst;
        _zz_io_output_payload_write = io_inputs_1_payload_write;
      end
      default : begin
        _zz_io_output_payload_addr_1 = io_inputs_2_payload_addr;
        _zz_io_output_payload_id = io_inputs_2_payload_id;
        _zz_io_output_payload_len = io_inputs_2_payload_len;
        _zz_io_output_payload_size = io_inputs_2_payload_size;
        _zz_io_output_payload_burst = io_inputs_2_payload_burst;
        _zz_io_output_payload_write = io_inputs_2_payload_write;
      end
    endcase
  end

  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign maskRouted_2 = (locked ? maskLocked_2 : maskProposal_2);
  assign _zz_maskProposal_0 = {io_inputs_2_valid,{io_inputs_1_valid,io_inputs_0_valid}};
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[5 : 3] | _zz_maskProposal_0_2[2 : 0]);
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign maskProposal_1 = _zz_maskProposal_0_3[1];
  assign maskProposal_2 = _zz_maskProposal_0_3[2];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_valid = (((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1)) || (io_inputs_2_valid && maskRouted_2));
  assign _zz_io_output_payload_addr = {maskRouted_2,maskRouted_1};
  assign io_output_payload_addr = _zz_io_output_payload_addr_1;
  assign io_output_payload_id = _zz_io_output_payload_id;
  assign io_output_payload_len = _zz_io_output_payload_len;
  assign io_output_payload_size = _zz_io_output_payload_size;
  assign io_output_payload_burst = _zz_io_output_payload_burst;
  assign io_output_payload_write = _zz_io_output_payload_write;
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_inputs_2_ready = (maskRouted_2 && io_output_ready);
  assign io_chosenOH = {maskRouted_2,{maskRouted_1,maskRouted_0}};
  assign _zz_io_chosen = io_chosenOH[1];
  assign _zz_io_chosen_1 = io_chosenOH[2];
  assign io_chosen = {_zz_io_chosen_1,_zz_io_chosen};
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b0;
      maskLocked_1 <= 1'b0;
      maskLocked_2 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
        maskLocked_2 <= maskRouted_2;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

module Axi4WriteOnlyErrorSlave_1 (
  input               io_axi_aw_valid,
  output              io_axi_aw_ready,
  input      [63:0]   io_axi_aw_payload_addr,
  input      [1:0]    io_axi_aw_payload_id,
  input      [7:0]    io_axi_aw_payload_len,
  input      [2:0]    io_axi_aw_payload_size,
  input      [1:0]    io_axi_aw_payload_burst,
  input               io_axi_w_valid,
  output              io_axi_w_ready,
  input      [63:0]   io_axi_w_payload_data,
  input      [7:0]    io_axi_w_payload_strb,
  input               io_axi_w_payload_last,
  output              io_axi_b_valid,
  input               io_axi_b_ready,
  output     [1:0]    io_axi_b_payload_id,
  output     [1:0]    io_axi_b_payload_resp,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  reg                 consumeData;
  reg                 sendRsp;
  reg        [1:0]    id;
  wire                io_axi_aw_fire;
  wire                io_axi_w_fire;
  wire                when_Axi4ErrorSlave_l24;
  wire                io_axi_b_fire;

  assign io_axi_aw_ready = (! (consumeData || sendRsp));
  assign io_axi_aw_fire = (io_axi_aw_valid && io_axi_aw_ready);
  assign io_axi_w_ready = consumeData;
  assign io_axi_w_fire = (io_axi_w_valid && io_axi_w_ready);
  assign when_Axi4ErrorSlave_l24 = (io_axi_w_fire && io_axi_w_payload_last);
  assign io_axi_b_valid = sendRsp;
  assign io_axi_b_payload_resp = 2'b11;
  assign io_axi_b_payload_id = id;
  assign io_axi_b_fire = (io_axi_b_valid && io_axi_b_ready);
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      consumeData <= 1'b0;
      sendRsp <= 1'b0;
    end else begin
      if(io_axi_aw_fire) begin
        consumeData <= 1'b1;
      end
      if(when_Axi4ErrorSlave_l24) begin
        consumeData <= 1'b0;
        sendRsp <= 1'b1;
      end
      if(io_axi_b_fire) begin
        sendRsp <= 1'b0;
      end
    end
  end

  always @(posedge io_axiClk) begin
    if(io_axi_aw_fire) begin
      id <= io_axi_aw_payload_id;
    end
  end


endmodule

//Axi4ReadOnlyErrorSlave_1 replaced by Axi4ReadOnlyErrorSlave_2

module Axi4ReadOnlyErrorSlave_2 (
  input               io_axi_ar_valid,
  output              io_axi_ar_ready,
  input      [63:0]   io_axi_ar_payload_addr,
  input      [1:0]    io_axi_ar_payload_id,
  input      [7:0]    io_axi_ar_payload_len,
  input      [2:0]    io_axi_ar_payload_size,
  input      [1:0]    io_axi_ar_payload_burst,
  output              io_axi_r_valid,
  input               io_axi_r_ready,
  output     [63:0]   io_axi_r_payload_data,
  output     [1:0]    io_axi_r_payload_id,
  output     [1:0]    io_axi_r_payload_resp,
  output              io_axi_r_payload_last,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  reg                 sendRsp;
  reg        [1:0]    id;
  reg        [7:0]    remaining;
  wire                remainingZero;
  wire                io_axi_ar_fire;

  assign remainingZero = (remaining == 8'h0);
  assign io_axi_ar_ready = (! sendRsp);
  assign io_axi_ar_fire = (io_axi_ar_valid && io_axi_ar_ready);
  assign io_axi_r_valid = sendRsp;
  assign io_axi_r_payload_id = id;
  assign io_axi_r_payload_resp = 2'b11;
  assign io_axi_r_payload_last = remainingZero;
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      sendRsp <= 1'b0;
    end else begin
      if(io_axi_ar_fire) begin
        sendRsp <= 1'b1;
      end
      if(sendRsp) begin
        if(io_axi_r_ready) begin
          if(remainingZero) begin
            sendRsp <= 1'b0;
          end
        end
      end
    end
  end

  always @(posedge io_axiClk) begin
    if(io_axi_ar_fire) begin
      remaining <= io_axi_ar_payload_len;
      id <= io_axi_ar_payload_id;
    end
    if(sendRsp) begin
      if(io_axi_r_ready) begin
        remaining <= (remaining - 8'h01);
      end
    end
  end


endmodule

module Axi4WriteOnlyDownsizer (
  input               io_input_aw_valid,
  output              io_input_aw_ready,
  input      [31:0]   io_input_aw_payload_addr,
  input      [3:0]    io_input_aw_payload_id,
  input      [3:0]    io_input_aw_payload_region,
  input      [7:0]    io_input_aw_payload_len,
  input      [2:0]    io_input_aw_payload_size,
  input      [1:0]    io_input_aw_payload_burst,
  input      [0:0]    io_input_aw_payload_lock,
  input      [3:0]    io_input_aw_payload_cache,
  input      [3:0]    io_input_aw_payload_qos,
  input      [2:0]    io_input_aw_payload_prot,
  input               io_input_w_valid,
  output              io_input_w_ready,
  input      [63:0]   io_input_w_payload_data,
  input      [7:0]    io_input_w_payload_strb,
  input               io_input_w_payload_last,
  output              io_input_b_valid,
  input               io_input_b_ready,
  output     [3:0]    io_input_b_payload_id,
  output     [1:0]    io_input_b_payload_resp,
  output              io_output_aw_valid,
  input               io_output_aw_ready,
  output     [31:0]   io_output_aw_payload_addr,
  output     [3:0]    io_output_aw_payload_id,
  output     [3:0]    io_output_aw_payload_region,
  output     [7:0]    io_output_aw_payload_len,
  output     [2:0]    io_output_aw_payload_size,
  output     [1:0]    io_output_aw_payload_burst,
  output     [0:0]    io_output_aw_payload_lock,
  output     [3:0]    io_output_aw_payload_cache,
  output     [3:0]    io_output_aw_payload_qos,
  output     [2:0]    io_output_aw_payload_prot,
  output              io_output_w_valid,
  input               io_output_w_ready,
  output     [31:0]   io_output_w_payload_data,
  output     [3:0]    io_output_w_payload_strb,
  output              io_output_w_payload_last,
  input               io_output_b_valid,
  output              io_output_b_ready,
  input      [3:0]    io_output_b_payload_id,
  input      [1:0]    io_output_b_payload_resp,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  wire                generator_io_input_ready;
  wire                generator_io_output_valid;
  wire       [31:0]   generator_io_output_payload_addr;
  wire       [3:0]    generator_io_output_payload_id;
  wire       [3:0]    generator_io_output_payload_region;
  wire       [7:0]    generator_io_output_payload_len;
  wire       [2:0]    generator_io_output_payload_size;
  wire       [1:0]    generator_io_output_payload_burst;
  wire       [0:0]    generator_io_output_payload_lock;
  wire       [3:0]    generator_io_output_payload_cache;
  wire       [3:0]    generator_io_output_payload_qos;
  wire       [2:0]    generator_io_output_payload_prot;
  wire       [31:0]   generator_io_start;
  wire       [6:0]    generator_io_ratio;
  wire       [2:0]    generator_io_size;
  wire                generator_io_working;
  wire                generator_io_last;
  wire                generator_io_done;
  wire                inputDataCounter_io_available;
  wire                inputDataCounter_io_working;
  wire                inputDataCounter_io_last;
  wire                inputDataCounter_io_done;
  wire       [7:0]    inputDataCounter_io_value;
  wire                streamCounter_io_available;
  wire                streamCounter_io_working;
  wire                streamCounter_io_last;
  wire                streamCounter_io_done;
  wire       [7:0]    streamCounter_io_value;
  wire                dataExtender_io_input_ready;
  wire                dataExtender_io_output_valid;
  wire       [63:0]   dataExtender_io_output_payload_data;
  wire       [7:0]    dataExtender_io_output_payload_strb;
  wire                dataExtender_io_output_payload_last;
  wire                dataExtender_io_working;
  wire                dataExtender_io_first;
  wire                dataExtender_io_last;
  wire                dataExtender_io_done;
  wire                rspCtrlStream_fifo_io_push_ready;
  wire                rspCtrlStream_fifo_io_pop_valid;
  wire                rspCtrlStream_fifo_io_pop_payload;
  wire       [1:0]    rspCtrlStream_fifo_io_occupancy;
  wire       [1:0]    rspCtrlStream_fifo_io_availability;
  wire       [7:0]    _zz_beatOffsetReg;
  wire       [7:0]    _zz_beatOffsetReg_1;
  wire       [7:0]    _zz_beatOffsetReg_2;
  wire       [5:0]    _zz_writeStream_w_payload_data;
  wire                writeStream_aw_valid;
  wire                writeStream_aw_ready;
  wire       [31:0]   writeStream_aw_payload_addr;
  wire       [3:0]    writeStream_aw_payload_id;
  wire       [3:0]    writeStream_aw_payload_region;
  wire       [7:0]    writeStream_aw_payload_len;
  wire       [2:0]    writeStream_aw_payload_size;
  wire       [1:0]    writeStream_aw_payload_burst;
  wire       [0:0]    writeStream_aw_payload_lock;
  wire       [3:0]    writeStream_aw_payload_cache;
  wire       [3:0]    writeStream_aw_payload_qos;
  wire       [2:0]    writeStream_aw_payload_prot;
  wire                writeStream_w_valid;
  wire                writeStream_w_ready;
  wire       [31:0]   writeStream_w_payload_data;
  wire       [3:0]    writeStream_w_payload_strb;
  wire                writeStream_w_payload_last;
  wire                writeStream_b_valid;
  wire                writeStream_b_ready;
  wire       [3:0]    writeStream_b_payload_id;
  wire       [1:0]    writeStream_b_payload_resp;
  wire                dataWorking;
  wire                _zz_io_input_aw_ready;
  wire                writeCmd_valid;
  wire                writeCmd_ready;
  wire       [31:0]   writeCmd_payload_addr;
  wire       [3:0]    writeCmd_payload_id;
  wire       [3:0]    writeCmd_payload_region;
  wire       [7:0]    writeCmd_payload_len;
  wire       [2:0]    writeCmd_payload_size;
  wire       [1:0]    writeCmd_payload_burst;
  wire       [0:0]    writeCmd_payload_lock;
  wire       [3:0]    writeCmd_payload_cache;
  wire       [3:0]    writeCmd_payload_qos;
  wire       [2:0]    writeCmd_payload_prot;
  wire                cmdStream_valid;
  reg                 cmdStream_ready;
  wire       [31:0]   cmdStream_payload_addr;
  wire       [3:0]    cmdStream_payload_id;
  wire       [3:0]    cmdStream_payload_region;
  wire       [7:0]    cmdStream_payload_len;
  wire       [2:0]    cmdStream_payload_size;
  wire       [1:0]    cmdStream_payload_burst;
  wire       [0:0]    cmdStream_payload_lock;
  wire       [3:0]    cmdStream_payload_cache;
  wire       [3:0]    cmdStream_payload_qos;
  wire       [2:0]    cmdStream_payload_prot;
  wire                staleInputData;
  wire                _zz_io_input_w_ready;
  wire                writeData_valid;
  wire                writeData_ready;
  wire       [63:0]   writeData_payload_data;
  wire       [7:0]    writeData_payload_strb;
  wire                writeData_payload_last;
  wire                writeCmd_fire;
  wire                writeData_fire;
  wire                rspCountStream_valid;
  wire                rspCountStream_ready;
  wire       [31:0]   rspCountStream_payload_addr;
  wire       [3:0]    rspCountStream_payload_id;
  wire       [3:0]    rspCountStream_payload_region;
  wire       [7:0]    rspCountStream_payload_len;
  wire       [2:0]    rspCountStream_payload_size;
  wire       [1:0]    rspCountStream_payload_burst;
  wire       [0:0]    rspCountStream_payload_lock;
  wire       [3:0]    rspCountStream_payload_cache;
  wire       [3:0]    rspCountStream_payload_qos;
  wire       [2:0]    rspCountStream_payload_prot;
  wire                countCmdStream_valid;
  wire                countCmdStream_ready;
  wire       [31:0]   countCmdStream_payload_addr;
  wire       [3:0]    countCmdStream_payload_id;
  wire       [3:0]    countCmdStream_payload_region;
  wire       [7:0]    countCmdStream_payload_len;
  wire       [2:0]    countCmdStream_payload_size;
  wire       [1:0]    countCmdStream_payload_burst;
  wire       [0:0]    countCmdStream_payload_lock;
  wire       [3:0]    countCmdStream_payload_cache;
  wire       [3:0]    countCmdStream_payload_qos;
  wire       [2:0]    countCmdStream_payload_prot;
  wire                outCmdStream_valid;
  wire                outCmdStream_ready;
  wire       [31:0]   outCmdStream_payload_addr;
  wire       [3:0]    outCmdStream_payload_id;
  wire       [3:0]    outCmdStream_payload_region;
  wire       [7:0]    outCmdStream_payload_len;
  wire       [2:0]    outCmdStream_payload_size;
  wire       [1:0]    outCmdStream_payload_burst;
  wire       [0:0]    outCmdStream_payload_lock;
  wire       [3:0]    outCmdStream_payload_cache;
  wire       [3:0]    outCmdStream_payload_qos;
  wire       [2:0]    outCmdStream_payload_prot;
  reg                 cmdStream_fork3_logic_linkEnable_0;
  reg                 cmdStream_fork3_logic_linkEnable_1;
  reg                 cmdStream_fork3_logic_linkEnable_2;
  wire                when_Stream_l992;
  wire                when_Stream_l992_1;
  wire                when_Stream_l992_2;
  wire                rspCountStream_fire;
  wire                countCmdStream_fire;
  wire                outCmdStream_fire;
  wire                dataStream_valid;
  wire                dataStream_ready;
  wire       [63:0]   dataStream_payload_data;
  wire       [7:0]    dataStream_payload_strb;
  wire                dataStream_payload_last;
  wire                countCmdStream_fire_1;
  wire                dataStream_fire;
  wire                countCmdStream_fire_2;
  reg        [2:0]    beatOffsetReg;
  reg        [2:0]    beatOffset;
  wire                countCmdStream_fire_3;
  wire                dataStream_fire_1;
  wire       [2:0]    offset;
  wire                staleData;
  wire                _zz_writeStream_w_valid;
  wire                rspCtrlStream_valid;
  wire                rspCtrlStream_ready;
  wire                rspCtrlStream_payload;
  wire                rspStream_valid;
  reg                 rspStream_ready;
  wire                rspStream_payload_1;
  wire       [3:0]    rspStream_payload_2_id;
  wire       [1:0]    rspStream_payload_2_resp;
  wire                rspStream_fire;
  wire                rspStream_fire_1;
  wire                when_Stream_l438;
  reg                 rspStream_thrown_valid;
  wire                rspStream_thrown_ready;
  wire                rspStream_thrown_payload_1;
  wire       [3:0]    rspStream_thrown_payload_2_id;
  wire       [1:0]    rspStream_thrown_payload_2_resp;

  assign _zz_beatOffsetReg = (_zz_beatOffsetReg_1 + _zz_beatOffsetReg_2);
  assign _zz_beatOffsetReg_1 = {5'd0, beatOffset};
  assign _zz_beatOffsetReg_2 = ({7'd0,1'b1} <<< generator_io_size);
  assign _zz_writeStream_w_payload_data = ({3'd0,offset} <<< 3);
  Axi4DownsizerSubTransactionGenerator_1 generator (
    .io_input_valid           (writeCmd_valid                         ), //i
    .io_input_ready           (generator_io_input_ready               ), //o
    .io_input_payload_addr    (writeCmd_payload_addr[31:0]            ), //i
    .io_input_payload_id      (writeCmd_payload_id[3:0]               ), //i
    .io_input_payload_region  (writeCmd_payload_region[3:0]           ), //i
    .io_input_payload_len     (writeCmd_payload_len[7:0]              ), //i
    .io_input_payload_size    (writeCmd_payload_size[2:0]             ), //i
    .io_input_payload_burst   (writeCmd_payload_burst[1:0]            ), //i
    .io_input_payload_lock    (writeCmd_payload_lock                  ), //i
    .io_input_payload_cache   (writeCmd_payload_cache[3:0]            ), //i
    .io_input_payload_qos     (writeCmd_payload_qos[3:0]              ), //i
    .io_input_payload_prot    (writeCmd_payload_prot[2:0]             ), //i
    .io_output_valid          (generator_io_output_valid              ), //o
    .io_output_ready          (cmdStream_ready                        ), //i
    .io_output_payload_addr   (generator_io_output_payload_addr[31:0] ), //o
    .io_output_payload_id     (generator_io_output_payload_id[3:0]    ), //o
    .io_output_payload_region (generator_io_output_payload_region[3:0]), //o
    .io_output_payload_len    (generator_io_output_payload_len[7:0]   ), //o
    .io_output_payload_size   (generator_io_output_payload_size[2:0]  ), //o
    .io_output_payload_burst  (generator_io_output_payload_burst[1:0] ), //o
    .io_output_payload_lock   (generator_io_output_payload_lock       ), //o
    .io_output_payload_cache  (generator_io_output_payload_cache[3:0] ), //o
    .io_output_payload_qos    (generator_io_output_payload_qos[3:0]   ), //o
    .io_output_payload_prot   (generator_io_output_payload_prot[2:0]  ), //o
    .io_start                 (generator_io_start[31:0]               ), //o
    .io_ratio                 (generator_io_ratio[6:0]                ), //o
    .io_size                  (generator_io_size[2:0]                 ), //o
    .io_working               (generator_io_working                   ), //o
    .io_last                  (generator_io_last                      ), //o
    .io_done                  (generator_io_done                      ), //o
    .io_axiClk                (io_axiClk                              ), //i
    .resetCtrl_axiReset       (resetCtrl_axiReset                     )  //i
  );
  StreamTransactionCounter inputDataCounter (
    .io_ctrlFire        (writeCmd_fire                 ), //i
    .io_targetFire      (writeData_fire                ), //i
    .io_available       (inputDataCounter_io_available ), //o
    .io_count           (writeCmd_payload_len[7:0]     ), //i
    .io_working         (inputDataCounter_io_working   ), //o
    .io_last            (inputDataCounter_io_last      ), //o
    .io_done            (inputDataCounter_io_done      ), //o
    .io_value           (inputDataCounter_io_value[7:0]), //o
    .io_axiClk          (io_axiClk                     ), //i
    .resetCtrl_axiReset (resetCtrl_axiReset            )  //i
  );
  StreamTransactionCounter streamCounter (
    .io_ctrlFire        (countCmdStream_fire_1          ), //i
    .io_targetFire      (dataStream_fire                ), //i
    .io_available       (streamCounter_io_available     ), //o
    .io_count           (countCmdStream_payload_len[7:0]), //i
    .io_working         (streamCounter_io_working       ), //o
    .io_last            (streamCounter_io_last          ), //o
    .io_done            (streamCounter_io_done          ), //o
    .io_value           (streamCounter_io_value[7:0]    ), //o
    .io_axiClk          (io_axiClk                      ), //i
    .resetCtrl_axiReset (resetCtrl_axiReset             )  //i
  );
  StreamTransactionExtender dataExtender (
    .io_count               (generator_io_ratio[6:0]                  ), //i
    .io_input_valid         (writeData_valid                          ), //i
    .io_input_ready         (dataExtender_io_input_ready              ), //o
    .io_input_payload_data  (writeData_payload_data[63:0]             ), //i
    .io_input_payload_strb  (writeData_payload_strb[7:0]              ), //i
    .io_input_payload_last  (writeData_payload_last                   ), //i
    .io_output_valid        (dataExtender_io_output_valid             ), //o
    .io_output_ready        (dataStream_ready                         ), //i
    .io_output_payload_data (dataExtender_io_output_payload_data[63:0]), //o
    .io_output_payload_strb (dataExtender_io_output_payload_strb[7:0] ), //o
    .io_output_payload_last (dataExtender_io_output_payload_last      ), //o
    .io_working             (dataExtender_io_working                  ), //o
    .io_first               (dataExtender_io_first                    ), //o
    .io_last                (dataExtender_io_last                     ), //o
    .io_done                (dataExtender_io_done                     ), //o
    .io_axiClk              (io_axiClk                                ), //i
    .resetCtrl_axiReset     (resetCtrl_axiReset                       )  //i
  );
  StreamFifo rspCtrlStream_fifo (
    .io_push_valid      (rspCtrlStream_valid                    ), //i
    .io_push_ready      (rspCtrlStream_fifo_io_push_ready       ), //o
    .io_push_payload    (rspCtrlStream_payload                  ), //i
    .io_pop_valid       (rspCtrlStream_fifo_io_pop_valid        ), //o
    .io_pop_ready       (rspStream_fire                         ), //i
    .io_pop_payload     (rspCtrlStream_fifo_io_pop_payload      ), //o
    .io_flush           (1'b0                                   ), //i
    .io_occupancy       (rspCtrlStream_fifo_io_occupancy[1:0]   ), //o
    .io_availability    (rspCtrlStream_fifo_io_availability[1:0]), //o
    .io_axiClk          (io_axiClk                              ), //i
    .resetCtrl_axiReset (resetCtrl_axiReset                     )  //i
  );
  assign _zz_io_input_aw_ready = (! dataWorking);
  assign writeCmd_valid = (io_input_aw_valid && _zz_io_input_aw_ready);
  assign io_input_aw_ready = (writeCmd_ready && _zz_io_input_aw_ready);
  assign writeCmd_payload_addr = io_input_aw_payload_addr;
  assign writeCmd_payload_id = io_input_aw_payload_id;
  assign writeCmd_payload_region = io_input_aw_payload_region;
  assign writeCmd_payload_len = io_input_aw_payload_len;
  assign writeCmd_payload_size = io_input_aw_payload_size;
  assign writeCmd_payload_burst = io_input_aw_payload_burst;
  assign writeCmd_payload_lock = io_input_aw_payload_lock;
  assign writeCmd_payload_cache = io_input_aw_payload_cache;
  assign writeCmd_payload_qos = io_input_aw_payload_qos;
  assign writeCmd_payload_prot = io_input_aw_payload_prot;
  assign writeCmd_ready = generator_io_input_ready;
  assign cmdStream_valid = generator_io_output_valid;
  assign cmdStream_payload_addr = generator_io_output_payload_addr;
  assign cmdStream_payload_id = generator_io_output_payload_id;
  assign cmdStream_payload_region = generator_io_output_payload_region;
  assign cmdStream_payload_len = generator_io_output_payload_len;
  assign cmdStream_payload_size = generator_io_output_payload_size;
  assign cmdStream_payload_burst = generator_io_output_payload_burst;
  assign cmdStream_payload_lock = generator_io_output_payload_lock;
  assign cmdStream_payload_cache = generator_io_output_payload_cache;
  assign cmdStream_payload_qos = generator_io_output_payload_qos;
  assign cmdStream_payload_prot = generator_io_output_payload_prot;
  assign _zz_io_input_w_ready = (! staleInputData);
  assign writeData_valid = (io_input_w_valid && _zz_io_input_w_ready);
  assign io_input_w_ready = (writeData_ready && _zz_io_input_w_ready);
  assign writeData_payload_data = io_input_w_payload_data;
  assign writeData_payload_strb = io_input_w_payload_strb;
  assign writeData_payload_last = io_input_w_payload_last;
  assign writeCmd_fire = (writeCmd_valid && writeCmd_ready);
  assign writeData_fire = (writeData_valid && writeData_ready);
  assign staleInputData = (! inputDataCounter_io_working);
  always @(*) begin
    cmdStream_ready = 1'b1;
    if(when_Stream_l992) begin
      cmdStream_ready = 1'b0;
    end
    if(when_Stream_l992_1) begin
      cmdStream_ready = 1'b0;
    end
    if(when_Stream_l992_2) begin
      cmdStream_ready = 1'b0;
    end
  end

  assign when_Stream_l992 = ((! rspCountStream_ready) && cmdStream_fork3_logic_linkEnable_0);
  assign when_Stream_l992_1 = ((! countCmdStream_ready) && cmdStream_fork3_logic_linkEnable_1);
  assign when_Stream_l992_2 = ((! outCmdStream_ready) && cmdStream_fork3_logic_linkEnable_2);
  assign rspCountStream_valid = (cmdStream_valid && cmdStream_fork3_logic_linkEnable_0);
  assign rspCountStream_payload_addr = cmdStream_payload_addr;
  assign rspCountStream_payload_id = cmdStream_payload_id;
  assign rspCountStream_payload_region = cmdStream_payload_region;
  assign rspCountStream_payload_len = cmdStream_payload_len;
  assign rspCountStream_payload_size = cmdStream_payload_size;
  assign rspCountStream_payload_burst = cmdStream_payload_burst;
  assign rspCountStream_payload_lock = cmdStream_payload_lock;
  assign rspCountStream_payload_cache = cmdStream_payload_cache;
  assign rspCountStream_payload_qos = cmdStream_payload_qos;
  assign rspCountStream_payload_prot = cmdStream_payload_prot;
  assign rspCountStream_fire = (rspCountStream_valid && rspCountStream_ready);
  assign countCmdStream_valid = (cmdStream_valid && cmdStream_fork3_logic_linkEnable_1);
  assign countCmdStream_payload_addr = cmdStream_payload_addr;
  assign countCmdStream_payload_id = cmdStream_payload_id;
  assign countCmdStream_payload_region = cmdStream_payload_region;
  assign countCmdStream_payload_len = cmdStream_payload_len;
  assign countCmdStream_payload_size = cmdStream_payload_size;
  assign countCmdStream_payload_burst = cmdStream_payload_burst;
  assign countCmdStream_payload_lock = cmdStream_payload_lock;
  assign countCmdStream_payload_cache = cmdStream_payload_cache;
  assign countCmdStream_payload_qos = cmdStream_payload_qos;
  assign countCmdStream_payload_prot = cmdStream_payload_prot;
  assign countCmdStream_fire = (countCmdStream_valid && countCmdStream_ready);
  assign outCmdStream_valid = (cmdStream_valid && cmdStream_fork3_logic_linkEnable_2);
  assign outCmdStream_payload_addr = cmdStream_payload_addr;
  assign outCmdStream_payload_id = cmdStream_payload_id;
  assign outCmdStream_payload_region = cmdStream_payload_region;
  assign outCmdStream_payload_len = cmdStream_payload_len;
  assign outCmdStream_payload_size = cmdStream_payload_size;
  assign outCmdStream_payload_burst = cmdStream_payload_burst;
  assign outCmdStream_payload_lock = cmdStream_payload_lock;
  assign outCmdStream_payload_cache = cmdStream_payload_cache;
  assign outCmdStream_payload_qos = cmdStream_payload_qos;
  assign outCmdStream_payload_prot = cmdStream_payload_prot;
  assign outCmdStream_fire = (outCmdStream_valid && outCmdStream_ready);
  assign writeStream_aw_valid = outCmdStream_valid;
  assign outCmdStream_ready = writeStream_aw_ready;
  assign writeStream_aw_payload_addr = outCmdStream_payload_addr;
  assign writeStream_aw_payload_id = outCmdStream_payload_id;
  assign writeStream_aw_payload_region = outCmdStream_payload_region;
  assign writeStream_aw_payload_len = outCmdStream_payload_len;
  assign writeStream_aw_payload_size = outCmdStream_payload_size;
  assign writeStream_aw_payload_burst = outCmdStream_payload_burst;
  assign writeStream_aw_payload_lock = outCmdStream_payload_lock;
  assign writeStream_aw_payload_cache = outCmdStream_payload_cache;
  assign writeStream_aw_payload_qos = outCmdStream_payload_qos;
  assign writeStream_aw_payload_prot = outCmdStream_payload_prot;
  assign countCmdStream_fire_1 = (countCmdStream_valid && countCmdStream_ready);
  assign dataStream_fire = (dataStream_valid && dataStream_ready);
  assign countCmdStream_ready = streamCounter_io_available;
  assign countCmdStream_fire_2 = (countCmdStream_valid && countCmdStream_ready);
  always @(*) begin
    beatOffset = beatOffsetReg;
    if(countCmdStream_fire_3) begin
      beatOffset = countCmdStream_payload_addr[2 : 0];
    end
  end

  assign countCmdStream_fire_3 = (countCmdStream_valid && countCmdStream_ready);
  assign dataStream_fire_1 = (dataStream_valid && dataStream_ready);
  assign offset = (beatOffset & (~ 3'b011));
  assign writeData_ready = dataExtender_io_input_ready;
  assign dataStream_valid = dataExtender_io_output_valid;
  assign dataStream_payload_data = dataExtender_io_output_payload_data;
  assign dataStream_payload_strb = dataExtender_io_output_payload_strb;
  assign dataStream_payload_last = dataExtender_io_output_payload_last;
  assign dataWorking = ((! inputDataCounter_io_available) || (! writeData_ready));
  assign staleData = (! streamCounter_io_working);
  assign _zz_writeStream_w_valid = (! staleData);
  assign dataStream_ready = (writeStream_w_ready && _zz_writeStream_w_valid);
  assign writeStream_w_valid = (dataStream_valid && _zz_writeStream_w_valid);
  assign writeStream_w_payload_data = dataStream_payload_data[_zz_writeStream_w_payload_data +: 32];
  assign writeStream_w_payload_last = streamCounter_io_last;
  assign writeStream_w_payload_strb = dataStream_payload_strb[offset +: 4];
  assign rspCtrlStream_valid = rspCountStream_valid;
  assign rspCountStream_ready = rspCtrlStream_ready;
  assign rspCtrlStream_payload = generator_io_last;
  assign rspCtrlStream_ready = rspCtrlStream_fifo_io_push_ready;
  assign rspStream_valid = (rspCtrlStream_fifo_io_pop_valid && writeStream_b_valid);
  assign rspStream_fire = (rspStream_valid && rspStream_ready);
  assign rspStream_fire_1 = (rspStream_valid && rspStream_ready);
  assign writeStream_b_ready = rspStream_fire_1;
  assign rspStream_payload_1 = rspCtrlStream_fifo_io_pop_payload;
  assign rspStream_payload_2_id = writeStream_b_payload_id;
  assign rspStream_payload_2_resp = writeStream_b_payload_resp;
  assign when_Stream_l438 = (! rspStream_payload_1);
  always @(*) begin
    rspStream_thrown_valid = rspStream_valid;
    if(when_Stream_l438) begin
      rspStream_thrown_valid = 1'b0;
    end
  end

  always @(*) begin
    rspStream_ready = rspStream_thrown_ready;
    if(when_Stream_l438) begin
      rspStream_ready = 1'b1;
    end
  end

  assign rspStream_thrown_payload_2_id = rspStream_payload_2_id;
  assign rspStream_thrown_payload_2_resp = rspStream_payload_2_resp;
  assign rspStream_thrown_payload_1 = rspStream_payload_1;
  assign io_input_b_valid = rspStream_thrown_valid;
  assign rspStream_thrown_ready = io_input_b_ready;
  assign io_input_b_payload_id = rspStream_thrown_payload_2_id;
  assign io_input_b_payload_resp = rspStream_thrown_payload_2_resp;
  assign io_output_aw_valid = writeStream_aw_valid;
  assign writeStream_aw_ready = io_output_aw_ready;
  assign io_output_aw_payload_addr = writeStream_aw_payload_addr;
  assign io_output_aw_payload_id = writeStream_aw_payload_id;
  assign io_output_aw_payload_region = writeStream_aw_payload_region;
  assign io_output_aw_payload_len = writeStream_aw_payload_len;
  assign io_output_aw_payload_size = writeStream_aw_payload_size;
  assign io_output_aw_payload_burst = writeStream_aw_payload_burst;
  assign io_output_aw_payload_lock = writeStream_aw_payload_lock;
  assign io_output_aw_payload_cache = writeStream_aw_payload_cache;
  assign io_output_aw_payload_qos = writeStream_aw_payload_qos;
  assign io_output_aw_payload_prot = writeStream_aw_payload_prot;
  assign io_output_w_valid = writeStream_w_valid;
  assign writeStream_w_ready = io_output_w_ready;
  assign io_output_w_payload_data = writeStream_w_payload_data;
  assign io_output_w_payload_strb = writeStream_w_payload_strb;
  assign io_output_w_payload_last = writeStream_w_payload_last;
  assign writeStream_b_valid = io_output_b_valid;
  assign io_output_b_ready = writeStream_b_ready;
  assign writeStream_b_payload_id = io_output_b_payload_id;
  assign writeStream_b_payload_resp = io_output_b_payload_resp;
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      cmdStream_fork3_logic_linkEnable_0 <= 1'b1;
      cmdStream_fork3_logic_linkEnable_1 <= 1'b1;
      cmdStream_fork3_logic_linkEnable_2 <= 1'b1;
    end else begin
      if(rspCountStream_fire) begin
        cmdStream_fork3_logic_linkEnable_0 <= 1'b0;
      end
      if(countCmdStream_fire) begin
        cmdStream_fork3_logic_linkEnable_1 <= 1'b0;
      end
      if(outCmdStream_fire) begin
        cmdStream_fork3_logic_linkEnable_2 <= 1'b0;
      end
      if(cmdStream_ready) begin
        cmdStream_fork3_logic_linkEnable_0 <= 1'b1;
        cmdStream_fork3_logic_linkEnable_1 <= 1'b1;
        cmdStream_fork3_logic_linkEnable_2 <= 1'b1;
      end
    end
  end

  always @(posedge io_axiClk) begin
    if(countCmdStream_fire_2) begin
      beatOffsetReg <= countCmdStream_payload_addr[2 : 0];
    end
    if(dataStream_fire_1) begin
      beatOffsetReg <= _zz_beatOffsetReg[2:0];
    end
  end


endmodule

module Axi4ReadOnlyDownsizer (
  input               io_input_ar_valid,
  output              io_input_ar_ready,
  input      [31:0]   io_input_ar_payload_addr,
  input      [3:0]    io_input_ar_payload_id,
  input      [3:0]    io_input_ar_payload_region,
  input      [7:0]    io_input_ar_payload_len,
  input      [2:0]    io_input_ar_payload_size,
  input      [1:0]    io_input_ar_payload_burst,
  input      [0:0]    io_input_ar_payload_lock,
  input      [3:0]    io_input_ar_payload_cache,
  input      [3:0]    io_input_ar_payload_qos,
  input      [2:0]    io_input_ar_payload_prot,
  output              io_input_r_valid,
  input               io_input_r_ready,
  output     [63:0]   io_input_r_payload_data,
  output     [3:0]    io_input_r_payload_id,
  output     [1:0]    io_input_r_payload_resp,
  output              io_input_r_payload_last,
  output              io_output_ar_valid,
  input               io_output_ar_ready,
  output     [31:0]   io_output_ar_payload_addr,
  output     [3:0]    io_output_ar_payload_id,
  output     [3:0]    io_output_ar_payload_region,
  output     [7:0]    io_output_ar_payload_len,
  output     [2:0]    io_output_ar_payload_size,
  output     [1:0]    io_output_ar_payload_burst,
  output     [0:0]    io_output_ar_payload_lock,
  output     [3:0]    io_output_ar_payload_cache,
  output     [3:0]    io_output_ar_payload_qos,
  output     [2:0]    io_output_ar_payload_prot,
  input               io_output_r_valid,
  output reg          io_output_r_ready,
  input      [31:0]   io_output_r_payload_data,
  input      [3:0]    io_output_r_payload_id,
  input      [1:0]    io_output_r_payload_resp,
  input               io_output_r_payload_last,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  wire                generator_io_input_ready;
  wire                generator_io_output_valid;
  wire       [31:0]   generator_io_output_payload_addr;
  wire       [3:0]    generator_io_output_payload_id;
  wire       [3:0]    generator_io_output_payload_region;
  wire       [7:0]    generator_io_output_payload_len;
  wire       [2:0]    generator_io_output_payload_size;
  wire       [1:0]    generator_io_output_payload_burst;
  wire       [0:0]    generator_io_output_payload_lock;
  wire       [3:0]    generator_io_output_payload_cache;
  wire       [3:0]    generator_io_output_payload_qos;
  wire       [2:0]    generator_io_output_payload_prot;
  wire       [31:0]   generator_io_start;
  wire       [6:0]    generator_io_ratio;
  wire       [2:0]    generator_io_size;
  wire                generator_io_working;
  wire                generator_io_last;
  wire                generator_io_done;
  wire                dataOutCounter_io_input_ready;
  wire                dataOutCounter_io_output_valid;
  wire       [6:0]    dataOutCounter_io_output_payload_ratio;
  wire       [2:0]    dataOutCounter_io_output_payload_size;
  wire       [7:0]    dataOutCounter_io_output_payload_len;
  wire       [31:0]   dataOutCounter_io_output_payload_start;
  wire                dataOutCounter_io_working;
  wire                dataOutCounter_io_first;
  wire                dataOutCounter_io_last;
  wire                dataOutCounter_io_done;
  wire                dataCounter_io_input_ready;
  wire                dataCounter_io_output_valid;
  wire       [6:0]    dataCounter_io_output_payload_ratio;
  wire       [2:0]    dataCounter_io_output_payload_size;
  wire       [7:0]    dataCounter_io_output_payload_len;
  wire       [31:0]   dataCounter_io_output_payload_start;
  wire                dataCounter_io_working;
  wire                dataCounter_io_first;
  wire                dataCounter_io_last;
  wire                dataCounter_io_done;
  wire       [7:0]    _zz_beatOffset;
  wire       [7:0]    _zz_beatOffset_1;
  wire       [7:0]    _zz_beatOffset_2;
  wire       [5:0]    _zz_dataReg_aheadValue;
  (* nowrshmsk *) reg        [63:0]   dataReg_aheadValue;
  wire                readCmdGen_valid;
  wire                readCmdGen_ready;
  wire       [31:0]   readCmdGen_payload_addr;
  wire       [3:0]    readCmdGen_payload_id;
  wire       [3:0]    readCmdGen_payload_region;
  wire       [7:0]    readCmdGen_payload_len;
  wire       [2:0]    readCmdGen_payload_size;
  wire       [1:0]    readCmdGen_payload_burst;
  wire       [0:0]    readCmdGen_payload_lock;
  wire       [3:0]    readCmdGen_payload_cache;
  wire       [3:0]    readCmdGen_payload_qos;
  wire       [2:0]    readCmdGen_payload_prot;
  wire                readCmdCount_valid;
  wire                readCmdCount_ready;
  wire       [31:0]   readCmdCount_payload_addr;
  wire       [3:0]    readCmdCount_payload_id;
  wire       [3:0]    readCmdCount_payload_region;
  wire       [7:0]    readCmdCount_payload_len;
  wire       [2:0]    readCmdCount_payload_size;
  wire       [1:0]    readCmdCount_payload_burst;
  wire       [0:0]    readCmdCount_payload_lock;
  wire       [3:0]    readCmdCount_payload_cache;
  wire       [3:0]    readCmdCount_payload_qos;
  wire       [2:0]    readCmdCount_payload_prot;
  wire                cmdStream_valid;
  wire                cmdStream_ready;
  wire       [31:0]   cmdStream_payload_addr;
  wire       [3:0]    cmdStream_payload_id;
  wire       [3:0]    cmdStream_payload_region;
  wire       [7:0]    cmdStream_payload_len;
  wire       [2:0]    cmdStream_payload_size;
  wire       [1:0]    cmdStream_payload_burst;
  wire       [0:0]    cmdStream_payload_lock;
  wire       [3:0]    cmdStream_payload_cache;
  wire       [3:0]    cmdStream_payload_qos;
  wire       [2:0]    cmdStream_payload_prot;
  wire       [6:0]    cmdState_ratio;
  wire       [2:0]    cmdState_size;
  wire       [7:0]    cmdState_len;
  wire       [31:0]   cmdState_start;
  wire                countCmdStream_valid;
  wire                countCmdStream_ready;
  wire       [6:0]    countCmdStream_payload_ratio;
  wire       [2:0]    countCmdStream_payload_size;
  wire       [7:0]    countCmdStream_payload_len;
  wire       [31:0]   countCmdStream_payload_start;
  wire                countOutStream_valid;
  wire                countOutStream_ready;
  wire       [6:0]    countOutStream_payload_ratio;
  wire       [2:0]    countOutStream_payload_size;
  wire       [7:0]    countOutStream_payload_len;
  wire       [31:0]   countOutStream_payload_start;
  wire                countStream_valid;
  wire                countStream_ready;
  wire       [6:0]    countStream_payload_ratio;
  wire       [2:0]    countStream_payload_size;
  wire       [7:0]    countStream_payload_len;
  wire       [31:0]   countStream_payload_start;
  wire                io_output_r_fire;
  reg        [63:0]   dataReg;
  reg        [2:0]    beatOffset;
  wire                countOutStream_fire;
  wire                when_Axi4Downsizer_l219;
  wire                io_output_r_fire_1;
  wire       [2:0]    offset;
  wire                dataOut_valid;
  wire                dataOut_ready;
  wire       [63:0]   dataOut_payload_data;
  wire       [3:0]    dataOut_payload_id;
  wire       [1:0]    dataOut_payload_resp;
  wire                dataOut_payload_last;
  reg                 lastLast;
  wire                countOutStream_fire_1;
  wire                when_Axi4Downsizer_l234;
  wire                io_output_r_fire_2;
  wire                when_Axi4Downsizer_l236;
  wire                when_Stream_l438;
  reg                 io_output_r_thrown_valid;
  wire                io_output_r_thrown_ready;
  wire       [31:0]   io_output_r_thrown_payload_data;
  wire       [3:0]    io_output_r_thrown_payload_id;
  wire       [1:0]    io_output_r_thrown_payload_resp;
  wire                io_output_r_thrown_payload_last;

  assign _zz_dataReg_aheadValue = ({3'd0,offset} <<< 3);
  assign _zz_beatOffset = (_zz_beatOffset_1 + _zz_beatOffset_2);
  assign _zz_beatOffset_1 = {5'd0, beatOffset};
  assign _zz_beatOffset_2 = ({7'd0,1'b1} <<< countStream_payload_size);
  Axi4DownsizerSubTransactionGenerator_1 generator (
    .io_input_valid           (readCmdGen_valid                       ), //i
    .io_input_ready           (generator_io_input_ready               ), //o
    .io_input_payload_addr    (readCmdGen_payload_addr[31:0]          ), //i
    .io_input_payload_id      (readCmdGen_payload_id[3:0]             ), //i
    .io_input_payload_region  (readCmdGen_payload_region[3:0]         ), //i
    .io_input_payload_len     (readCmdGen_payload_len[7:0]            ), //i
    .io_input_payload_size    (readCmdGen_payload_size[2:0]           ), //i
    .io_input_payload_burst   (readCmdGen_payload_burst[1:0]          ), //i
    .io_input_payload_lock    (readCmdGen_payload_lock                ), //i
    .io_input_payload_cache   (readCmdGen_payload_cache[3:0]          ), //i
    .io_input_payload_qos     (readCmdGen_payload_qos[3:0]            ), //i
    .io_input_payload_prot    (readCmdGen_payload_prot[2:0]           ), //i
    .io_output_valid          (generator_io_output_valid              ), //o
    .io_output_ready          (cmdStream_ready                        ), //i
    .io_output_payload_addr   (generator_io_output_payload_addr[31:0] ), //o
    .io_output_payload_id     (generator_io_output_payload_id[3:0]    ), //o
    .io_output_payload_region (generator_io_output_payload_region[3:0]), //o
    .io_output_payload_len    (generator_io_output_payload_len[7:0]   ), //o
    .io_output_payload_size   (generator_io_output_payload_size[2:0]  ), //o
    .io_output_payload_burst  (generator_io_output_payload_burst[1:0] ), //o
    .io_output_payload_lock   (generator_io_output_payload_lock       ), //o
    .io_output_payload_cache  (generator_io_output_payload_cache[3:0] ), //o
    .io_output_payload_qos    (generator_io_output_payload_qos[3:0]   ), //o
    .io_output_payload_prot   (generator_io_output_payload_prot[2:0]  ), //o
    .io_start                 (generator_io_start[31:0]               ), //o
    .io_ratio                 (generator_io_ratio[6:0]                ), //o
    .io_size                  (generator_io_size[2:0]                 ), //o
    .io_working               (generator_io_working                   ), //o
    .io_last                  (generator_io_last                      ), //o
    .io_done                  (generator_io_done                      ), //o
    .io_axiClk                (io_axiClk                              ), //i
    .resetCtrl_axiReset       (resetCtrl_axiReset                     )  //i
  );
  StreamTransactionExtender_1 dataOutCounter (
    .io_count                (countCmdStream_payload_len[7:0]             ), //i
    .io_input_valid          (countCmdStream_valid                        ), //i
    .io_input_ready          (dataOutCounter_io_input_ready               ), //o
    .io_input_payload_ratio  (countCmdStream_payload_ratio[6:0]           ), //i
    .io_input_payload_size   (countCmdStream_payload_size[2:0]            ), //i
    .io_input_payload_len    (countCmdStream_payload_len[7:0]             ), //i
    .io_input_payload_start  (countCmdStream_payload_start[31:0]          ), //i
    .io_output_valid         (dataOutCounter_io_output_valid              ), //o
    .io_output_ready         (countOutStream_ready                        ), //i
    .io_output_payload_ratio (dataOutCounter_io_output_payload_ratio[6:0] ), //o
    .io_output_payload_size  (dataOutCounter_io_output_payload_size[2:0]  ), //o
    .io_output_payload_len   (dataOutCounter_io_output_payload_len[7:0]   ), //o
    .io_output_payload_start (dataOutCounter_io_output_payload_start[31:0]), //o
    .io_working              (dataOutCounter_io_working                   ), //o
    .io_first                (dataOutCounter_io_first                     ), //o
    .io_last                 (dataOutCounter_io_last                      ), //o
    .io_done                 (dataOutCounter_io_done                      ), //o
    .io_axiClk               (io_axiClk                                   ), //i
    .resetCtrl_axiReset      (resetCtrl_axiReset                          )  //i
  );
  StreamTransactionExtender_2 dataCounter (
    .io_count                (countOutStream_payload_ratio[6:0]        ), //i
    .io_input_valid          (countOutStream_valid                     ), //i
    .io_input_ready          (dataCounter_io_input_ready               ), //o
    .io_input_payload_ratio  (countOutStream_payload_ratio[6:0]        ), //i
    .io_input_payload_size   (countOutStream_payload_size[2:0]         ), //i
    .io_input_payload_len    (countOutStream_payload_len[7:0]          ), //i
    .io_input_payload_start  (countOutStream_payload_start[31:0]       ), //i
    .io_output_valid         (dataCounter_io_output_valid              ), //o
    .io_output_ready         (countStream_ready                        ), //i
    .io_output_payload_ratio (dataCounter_io_output_payload_ratio[6:0] ), //o
    .io_output_payload_size  (dataCounter_io_output_payload_size[2:0]  ), //o
    .io_output_payload_len   (dataCounter_io_output_payload_len[7:0]   ), //o
    .io_output_payload_start (dataCounter_io_output_payload_start[31:0]), //o
    .io_working              (dataCounter_io_working                   ), //o
    .io_first                (dataCounter_io_first                     ), //o
    .io_last                 (dataCounter_io_last                      ), //o
    .io_done                 (dataCounter_io_done                      ), //o
    .io_axiClk               (io_axiClk                                ), //i
    .resetCtrl_axiReset      (resetCtrl_axiReset                       )  //i
  );
  always @(*) begin
    dataReg_aheadValue = dataReg;
    if(io_output_r_valid) begin
      dataReg_aheadValue[_zz_dataReg_aheadValue +: 32] = io_output_r_payload_data;
    end
  end

  assign io_input_ar_ready = (readCmdGen_ready && readCmdCount_ready);
  assign readCmdGen_valid = (io_input_ar_valid && io_input_ar_ready);
  assign readCmdCount_valid = (io_input_ar_valid && io_input_ar_ready);
  assign readCmdGen_payload_addr = io_input_ar_payload_addr;
  assign readCmdGen_payload_id = io_input_ar_payload_id;
  assign readCmdGen_payload_region = io_input_ar_payload_region;
  assign readCmdGen_payload_len = io_input_ar_payload_len;
  assign readCmdGen_payload_size = io_input_ar_payload_size;
  assign readCmdGen_payload_burst = io_input_ar_payload_burst;
  assign readCmdGen_payload_lock = io_input_ar_payload_lock;
  assign readCmdGen_payload_cache = io_input_ar_payload_cache;
  assign readCmdGen_payload_qos = io_input_ar_payload_qos;
  assign readCmdGen_payload_prot = io_input_ar_payload_prot;
  assign readCmdCount_payload_addr = io_input_ar_payload_addr;
  assign readCmdCount_payload_id = io_input_ar_payload_id;
  assign readCmdCount_payload_region = io_input_ar_payload_region;
  assign readCmdCount_payload_len = io_input_ar_payload_len;
  assign readCmdCount_payload_size = io_input_ar_payload_size;
  assign readCmdCount_payload_burst = io_input_ar_payload_burst;
  assign readCmdCount_payload_lock = io_input_ar_payload_lock;
  assign readCmdCount_payload_cache = io_input_ar_payload_cache;
  assign readCmdCount_payload_qos = io_input_ar_payload_qos;
  assign readCmdCount_payload_prot = io_input_ar_payload_prot;
  assign readCmdGen_ready = generator_io_input_ready;
  assign cmdStream_valid = generator_io_output_valid;
  assign cmdStream_payload_addr = generator_io_output_payload_addr;
  assign cmdStream_payload_id = generator_io_output_payload_id;
  assign cmdStream_payload_region = generator_io_output_payload_region;
  assign cmdStream_payload_len = generator_io_output_payload_len;
  assign cmdStream_payload_size = generator_io_output_payload_size;
  assign cmdStream_payload_burst = generator_io_output_payload_burst;
  assign cmdStream_payload_lock = generator_io_output_payload_lock;
  assign cmdStream_payload_cache = generator_io_output_payload_cache;
  assign cmdStream_payload_qos = generator_io_output_payload_qos;
  assign cmdStream_payload_prot = generator_io_output_payload_prot;
  assign io_output_ar_valid = cmdStream_valid;
  assign cmdStream_ready = io_output_ar_ready;
  assign io_output_ar_payload_addr = cmdStream_payload_addr;
  assign io_output_ar_payload_id = cmdStream_payload_id;
  assign io_output_ar_payload_region = cmdStream_payload_region;
  assign io_output_ar_payload_len = cmdStream_payload_len;
  assign io_output_ar_payload_size = cmdStream_payload_size;
  assign io_output_ar_payload_burst = cmdStream_payload_burst;
  assign io_output_ar_payload_lock = cmdStream_payload_lock;
  assign io_output_ar_payload_cache = cmdStream_payload_cache;
  assign io_output_ar_payload_qos = cmdStream_payload_qos;
  assign io_output_ar_payload_prot = cmdStream_payload_prot;
  assign countCmdStream_valid = readCmdCount_valid;
  assign readCmdCount_ready = countCmdStream_ready;
  assign countCmdStream_payload_ratio = generator_io_ratio;
  assign countCmdStream_payload_size = generator_io_size;
  assign countCmdStream_payload_len = readCmdCount_payload_len;
  assign countCmdStream_payload_start = generator_io_start;
  assign countCmdStream_ready = dataOutCounter_io_input_ready;
  assign countOutStream_valid = dataOutCounter_io_output_valid;
  assign countOutStream_payload_ratio = dataOutCounter_io_output_payload_ratio;
  assign countOutStream_payload_size = dataOutCounter_io_output_payload_size;
  assign countOutStream_payload_len = dataOutCounter_io_output_payload_len;
  assign countOutStream_payload_start = dataOutCounter_io_output_payload_start;
  assign countOutStream_ready = dataCounter_io_input_ready;
  assign countStream_valid = dataCounter_io_output_valid;
  assign countStream_payload_ratio = dataCounter_io_output_payload_ratio;
  assign countStream_payload_size = dataCounter_io_output_payload_size;
  assign countStream_payload_len = dataCounter_io_output_payload_len;
  assign countStream_payload_start = dataCounter_io_output_payload_start;
  assign io_output_r_fire = (io_output_r_valid && io_output_r_ready);
  assign countStream_ready = io_output_r_fire;
  assign countOutStream_fire = (countOutStream_valid && countOutStream_ready);
  assign when_Axi4Downsizer_l219 = (countOutStream_fire && dataOutCounter_io_first);
  assign io_output_r_fire_1 = (io_output_r_valid && io_output_r_ready);
  assign offset = (beatOffset & (~ 3'b011));
  assign countOutStream_fire_1 = (countOutStream_valid && countOutStream_ready);
  assign when_Axi4Downsizer_l234 = ((dataOutCounter_io_working && dataOutCounter_io_last) && countOutStream_fire_1);
  assign io_output_r_fire_2 = (io_output_r_valid && io_output_r_ready);
  assign when_Axi4Downsizer_l236 = (dataCounter_io_last && io_output_r_fire_2);
  assign when_Stream_l438 = (! dataCounter_io_last);
  always @(*) begin
    io_output_r_thrown_valid = io_output_r_valid;
    if(when_Stream_l438) begin
      io_output_r_thrown_valid = 1'b0;
    end
  end

  always @(*) begin
    io_output_r_ready = io_output_r_thrown_ready;
    if(when_Stream_l438) begin
      io_output_r_ready = 1'b1;
    end
  end

  assign io_output_r_thrown_payload_data = io_output_r_payload_data;
  assign io_output_r_thrown_payload_id = io_output_r_payload_id;
  assign io_output_r_thrown_payload_resp = io_output_r_payload_resp;
  assign io_output_r_thrown_payload_last = io_output_r_payload_last;
  assign dataOut_valid = io_output_r_thrown_valid;
  assign io_output_r_thrown_ready = dataOut_ready;
  assign dataOut_payload_data = dataReg_aheadValue;
  assign dataOut_payload_last = (io_output_r_thrown_payload_last && lastLast);
  assign dataOut_payload_id = io_output_r_thrown_payload_id;
  assign dataOut_payload_resp = io_output_r_thrown_payload_resp;
  assign io_input_r_valid = dataOut_valid;
  assign dataOut_ready = io_input_r_ready;
  assign io_input_r_payload_data = dataOut_payload_data;
  assign io_input_r_payload_id = dataOut_payload_id;
  assign io_input_r_payload_resp = dataOut_payload_resp;
  assign io_input_r_payload_last = dataOut_payload_last;
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      dataReg <= 64'h0;
      beatOffset <= 3'b000;
      lastLast <= 1'b0;
    end else begin
      if(when_Axi4Downsizer_l219) begin
        beatOffset <= countOutStream_payload_start[2 : 0];
      end else begin
        if(io_output_r_fire_1) begin
          beatOffset <= _zz_beatOffset[2:0];
        end
      end
      if(when_Axi4Downsizer_l234) begin
        lastLast <= 1'b1;
      end else begin
        if(when_Axi4Downsizer_l236) begin
          lastLast <= 1'b0;
        end
      end
      dataReg <= dataReg_aheadValue;
    end
  end


endmodule

module SramBanks_1 (
  input               sram_0_ports_cmd_valid,
  input      [1:0]    sram_0_ports_cmd_payload_addr,
  input      [7:0]    sram_0_ports_cmd_payload_wen,
  input      [511:0]  sram_0_ports_cmd_payload_wdata,
  input      [63:0]   sram_0_ports_cmd_payload_wstrb,
  output              sram_0_ports_rsp_valid,
  output reg [511:0]  sram_0_ports_rsp_payload_data,
  input               sram_1_ports_cmd_valid,
  input      [1:0]    sram_1_ports_cmd_payload_addr,
  input      [7:0]    sram_1_ports_cmd_payload_wen,
  input      [511:0]  sram_1_ports_cmd_payload_wdata,
  input      [63:0]   sram_1_ports_cmd_payload_wstrb,
  output              sram_1_ports_rsp_valid,
  output reg [511:0]  sram_1_ports_rsp_payload_data,
  input               sram_2_ports_cmd_valid,
  input      [1:0]    sram_2_ports_cmd_payload_addr,
  input      [7:0]    sram_2_ports_cmd_payload_wen,
  input      [511:0]  sram_2_ports_cmd_payload_wdata,
  input      [63:0]   sram_2_ports_cmd_payload_wstrb,
  output              sram_2_ports_rsp_valid,
  output reg [511:0]  sram_2_ports_rsp_payload_data,
  input               sram_3_ports_cmd_valid,
  input      [1:0]    sram_3_ports_cmd_payload_addr,
  input      [7:0]    sram_3_ports_cmd_payload_wen,
  input      [511:0]  sram_3_ports_cmd_payload_wdata,
  input      [63:0]   sram_3_ports_cmd_payload_wstrb,
  output              sram_3_ports_rsp_valid,
  output reg [511:0]  sram_3_ports_rsp_payload_data,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  wire       [63:0]   _zz_sram_0_banks_0_bank_port1;
  wire       [63:0]   _zz_sram_0_banks_1_bank_port1;
  wire       [63:0]   _zz_sram_0_banks_2_bank_port1;
  wire       [63:0]   _zz_sram_0_banks_3_bank_port1;
  wire       [63:0]   _zz_sram_0_banks_4_bank_port1;
  wire       [63:0]   _zz_sram_0_banks_5_bank_port1;
  wire       [63:0]   _zz_sram_0_banks_6_bank_port1;
  wire       [63:0]   _zz_sram_0_banks_7_bank_port1;
  wire       [63:0]   _zz_sram_1_banks_0_bank_port1;
  wire       [63:0]   _zz_sram_1_banks_1_bank_port1;
  wire       [63:0]   _zz_sram_1_banks_2_bank_port1;
  wire       [63:0]   _zz_sram_1_banks_3_bank_port1;
  wire       [63:0]   _zz_sram_1_banks_4_bank_port1;
  wire       [63:0]   _zz_sram_1_banks_5_bank_port1;
  wire       [63:0]   _zz_sram_1_banks_6_bank_port1;
  wire       [63:0]   _zz_sram_1_banks_7_bank_port1;
  wire       [63:0]   _zz_sram_2_banks_0_bank_port1;
  wire       [63:0]   _zz_sram_2_banks_1_bank_port1;
  wire       [63:0]   _zz_sram_2_banks_2_bank_port1;
  wire       [63:0]   _zz_sram_2_banks_3_bank_port1;
  wire       [63:0]   _zz_sram_2_banks_4_bank_port1;
  wire       [63:0]   _zz_sram_2_banks_5_bank_port1;
  wire       [63:0]   _zz_sram_2_banks_6_bank_port1;
  wire       [63:0]   _zz_sram_2_banks_7_bank_port1;
  wire       [63:0]   _zz_sram_3_banks_0_bank_port1;
  wire       [63:0]   _zz_sram_3_banks_1_bank_port1;
  wire       [63:0]   _zz_sram_3_banks_2_bank_port1;
  wire       [63:0]   _zz_sram_3_banks_3_bank_port1;
  wire       [63:0]   _zz_sram_3_banks_4_bank_port1;
  wire       [63:0]   _zz_sram_3_banks_5_bank_port1;
  wire       [63:0]   _zz_sram_3_banks_6_bank_port1;
  wire       [63:0]   _zz_sram_3_banks_7_bank_port1;
  wire       [63:0]   _zz_sram_0_banks_0_bank_port;
  wire       [7:0]    _zz_sram_0_banks_0_bank_port_1;
  wire                _zz_sram_0_banks_0_bank_port_2;
  wire       [63:0]   _zz_sram_0_banks_1_bank_port;
  wire       [7:0]    _zz_sram_0_banks_1_bank_port_1;
  wire                _zz_sram_0_banks_1_bank_port_2;
  wire       [63:0]   _zz_sram_0_banks_2_bank_port;
  wire       [7:0]    _zz_sram_0_banks_2_bank_port_1;
  wire                _zz_sram_0_banks_2_bank_port_2;
  wire       [63:0]   _zz_sram_0_banks_3_bank_port;
  wire       [7:0]    _zz_sram_0_banks_3_bank_port_1;
  wire                _zz_sram_0_banks_3_bank_port_2;
  wire       [63:0]   _zz_sram_0_banks_4_bank_port;
  wire       [7:0]    _zz_sram_0_banks_4_bank_port_1;
  wire                _zz_sram_0_banks_4_bank_port_2;
  wire       [63:0]   _zz_sram_0_banks_5_bank_port;
  wire       [7:0]    _zz_sram_0_banks_5_bank_port_1;
  wire                _zz_sram_0_banks_5_bank_port_2;
  wire       [63:0]   _zz_sram_0_banks_6_bank_port;
  wire       [7:0]    _zz_sram_0_banks_6_bank_port_1;
  wire                _zz_sram_0_banks_6_bank_port_2;
  wire       [63:0]   _zz_sram_0_banks_7_bank_port;
  wire       [7:0]    _zz_sram_0_banks_7_bank_port_1;
  wire                _zz_sram_0_banks_7_bank_port_2;
  wire       [63:0]   _zz_sram_1_banks_0_bank_port;
  wire       [7:0]    _zz_sram_1_banks_0_bank_port_1;
  wire                _zz_sram_1_banks_0_bank_port_2;
  wire       [63:0]   _zz_sram_1_banks_1_bank_port;
  wire       [7:0]    _zz_sram_1_banks_1_bank_port_1;
  wire                _zz_sram_1_banks_1_bank_port_2;
  wire       [63:0]   _zz_sram_1_banks_2_bank_port;
  wire       [7:0]    _zz_sram_1_banks_2_bank_port_1;
  wire                _zz_sram_1_banks_2_bank_port_2;
  wire       [63:0]   _zz_sram_1_banks_3_bank_port;
  wire       [7:0]    _zz_sram_1_banks_3_bank_port_1;
  wire                _zz_sram_1_banks_3_bank_port_2;
  wire       [63:0]   _zz_sram_1_banks_4_bank_port;
  wire       [7:0]    _zz_sram_1_banks_4_bank_port_1;
  wire                _zz_sram_1_banks_4_bank_port_2;
  wire       [63:0]   _zz_sram_1_banks_5_bank_port;
  wire       [7:0]    _zz_sram_1_banks_5_bank_port_1;
  wire                _zz_sram_1_banks_5_bank_port_2;
  wire       [63:0]   _zz_sram_1_banks_6_bank_port;
  wire       [7:0]    _zz_sram_1_banks_6_bank_port_1;
  wire                _zz_sram_1_banks_6_bank_port_2;
  wire       [63:0]   _zz_sram_1_banks_7_bank_port;
  wire       [7:0]    _zz_sram_1_banks_7_bank_port_1;
  wire                _zz_sram_1_banks_7_bank_port_2;
  wire       [63:0]   _zz_sram_2_banks_0_bank_port;
  wire       [7:0]    _zz_sram_2_banks_0_bank_port_1;
  wire                _zz_sram_2_banks_0_bank_port_2;
  wire       [63:0]   _zz_sram_2_banks_1_bank_port;
  wire       [7:0]    _zz_sram_2_banks_1_bank_port_1;
  wire                _zz_sram_2_banks_1_bank_port_2;
  wire       [63:0]   _zz_sram_2_banks_2_bank_port;
  wire       [7:0]    _zz_sram_2_banks_2_bank_port_1;
  wire                _zz_sram_2_banks_2_bank_port_2;
  wire       [63:0]   _zz_sram_2_banks_3_bank_port;
  wire       [7:0]    _zz_sram_2_banks_3_bank_port_1;
  wire                _zz_sram_2_banks_3_bank_port_2;
  wire       [63:0]   _zz_sram_2_banks_4_bank_port;
  wire       [7:0]    _zz_sram_2_banks_4_bank_port_1;
  wire                _zz_sram_2_banks_4_bank_port_2;
  wire       [63:0]   _zz_sram_2_banks_5_bank_port;
  wire       [7:0]    _zz_sram_2_banks_5_bank_port_1;
  wire                _zz_sram_2_banks_5_bank_port_2;
  wire       [63:0]   _zz_sram_2_banks_6_bank_port;
  wire       [7:0]    _zz_sram_2_banks_6_bank_port_1;
  wire                _zz_sram_2_banks_6_bank_port_2;
  wire       [63:0]   _zz_sram_2_banks_7_bank_port;
  wire       [7:0]    _zz_sram_2_banks_7_bank_port_1;
  wire                _zz_sram_2_banks_7_bank_port_2;
  wire       [63:0]   _zz_sram_3_banks_0_bank_port;
  wire       [7:0]    _zz_sram_3_banks_0_bank_port_1;
  wire                _zz_sram_3_banks_0_bank_port_2;
  wire       [63:0]   _zz_sram_3_banks_1_bank_port;
  wire       [7:0]    _zz_sram_3_banks_1_bank_port_1;
  wire                _zz_sram_3_banks_1_bank_port_2;
  wire       [63:0]   _zz_sram_3_banks_2_bank_port;
  wire       [7:0]    _zz_sram_3_banks_2_bank_port_1;
  wire                _zz_sram_3_banks_2_bank_port_2;
  wire       [63:0]   _zz_sram_3_banks_3_bank_port;
  wire       [7:0]    _zz_sram_3_banks_3_bank_port_1;
  wire                _zz_sram_3_banks_3_bank_port_2;
  wire       [63:0]   _zz_sram_3_banks_4_bank_port;
  wire       [7:0]    _zz_sram_3_banks_4_bank_port_1;
  wire                _zz_sram_3_banks_4_bank_port_2;
  wire       [63:0]   _zz_sram_3_banks_5_bank_port;
  wire       [7:0]    _zz_sram_3_banks_5_bank_port_1;
  wire                _zz_sram_3_banks_5_bank_port_2;
  wire       [63:0]   _zz_sram_3_banks_6_bank_port;
  wire       [7:0]    _zz_sram_3_banks_6_bank_port_1;
  wire                _zz_sram_3_banks_6_bank_port_2;
  wire       [63:0]   _zz_sram_3_banks_7_bank_port;
  wire       [7:0]    _zz_sram_3_banks_7_bank_port_1;
  wire                _zz_sram_3_banks_7_bank_port_2;
  reg                 _zz_sram_0_ports_rsp_valid;
  wire                when_SramBanks_l75;
  reg                 _zz_sram_1_ports_rsp_valid;
  wire                when_SramBanks_l75_1;
  reg                 _zz_sram_2_ports_rsp_valid;
  wire                when_SramBanks_l75_2;
  reg                 _zz_sram_3_ports_rsp_valid;
  wire                when_SramBanks_l75_3;
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_0_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_0_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_0_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_0_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_0_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_0_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_0_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_0_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_1_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_1_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_1_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_1_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_1_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_1_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_1_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_1_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_2_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_2_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_2_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_2_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_2_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_2_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_2_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_2_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_3_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_3_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_3_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_3_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_3_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_3_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_3_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_3_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_4_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_4_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_4_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_4_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_4_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_4_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_4_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_4_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_5_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_5_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_5_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_5_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_5_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_5_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_5_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_5_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_6_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_6_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_6_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_6_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_6_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_6_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_6_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_6_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_7_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_7_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_7_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_7_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_7_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_7_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_7_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_7_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_0_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_0_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_0_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_0_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_0_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_0_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_0_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_0_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_1_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_1_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_1_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_1_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_1_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_1_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_1_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_1_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_2_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_2_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_2_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_2_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_2_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_2_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_2_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_2_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_3_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_3_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_3_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_3_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_3_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_3_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_3_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_3_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_4_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_4_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_4_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_4_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_4_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_4_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_4_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_4_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_5_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_5_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_5_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_5_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_5_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_5_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_5_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_5_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_6_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_6_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_6_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_6_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_6_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_6_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_6_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_6_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_7_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_7_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_7_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_7_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_7_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_7_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_7_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_7_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_0_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_0_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_0_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_0_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_0_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_0_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_0_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_0_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_1_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_1_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_1_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_1_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_1_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_1_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_1_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_1_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_2_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_2_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_2_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_2_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_2_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_2_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_2_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_2_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_3_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_3_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_3_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_3_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_3_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_3_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_3_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_3_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_4_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_4_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_4_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_4_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_4_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_4_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_4_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_4_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_5_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_5_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_5_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_5_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_5_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_5_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_5_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_5_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_6_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_6_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_6_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_6_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_6_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_6_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_6_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_6_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_7_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_7_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_7_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_7_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_7_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_7_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_7_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_7_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_0_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_0_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_0_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_0_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_0_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_0_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_0_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_0_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_1_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_1_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_1_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_1_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_1_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_1_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_1_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_1_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_2_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_2_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_2_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_2_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_2_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_2_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_2_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_2_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_3_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_3_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_3_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_3_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_3_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_3_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_3_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_3_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_4_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_4_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_4_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_4_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_4_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_4_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_4_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_4_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_5_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_5_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_5_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_5_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_5_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_5_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_5_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_5_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_6_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_6_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_6_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_6_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_6_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_6_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_6_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_6_bank_symbol7 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_7_bank_symbol0 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_7_bank_symbol1 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_7_bank_symbol2 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_7_bank_symbol3 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_7_bank_symbol4 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_7_bank_symbol5 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_7_bank_symbol6 [0:3];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_7_bank_symbol7 [0:3];

  assign _zz_sram_0_banks_0_bank_port = sram_0_ports_cmd_payload_wdata[63 : 0];
  assign _zz_sram_0_banks_0_bank_port_1 = sram_0_ports_cmd_payload_wstrb[7 : 0];
  assign _zz_sram_0_banks_0_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[0]);
  assign _zz_sram_0_banks_1_bank_port = sram_0_ports_cmd_payload_wdata[127 : 64];
  assign _zz_sram_0_banks_1_bank_port_1 = sram_0_ports_cmd_payload_wstrb[15 : 8];
  assign _zz_sram_0_banks_1_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[1]);
  assign _zz_sram_0_banks_2_bank_port = sram_0_ports_cmd_payload_wdata[191 : 128];
  assign _zz_sram_0_banks_2_bank_port_1 = sram_0_ports_cmd_payload_wstrb[23 : 16];
  assign _zz_sram_0_banks_2_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[2]);
  assign _zz_sram_0_banks_3_bank_port = sram_0_ports_cmd_payload_wdata[255 : 192];
  assign _zz_sram_0_banks_3_bank_port_1 = sram_0_ports_cmd_payload_wstrb[31 : 24];
  assign _zz_sram_0_banks_3_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[3]);
  assign _zz_sram_0_banks_4_bank_port = sram_0_ports_cmd_payload_wdata[319 : 256];
  assign _zz_sram_0_banks_4_bank_port_1 = sram_0_ports_cmd_payload_wstrb[39 : 32];
  assign _zz_sram_0_banks_4_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[4]);
  assign _zz_sram_0_banks_5_bank_port = sram_0_ports_cmd_payload_wdata[383 : 320];
  assign _zz_sram_0_banks_5_bank_port_1 = sram_0_ports_cmd_payload_wstrb[47 : 40];
  assign _zz_sram_0_banks_5_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[5]);
  assign _zz_sram_0_banks_6_bank_port = sram_0_ports_cmd_payload_wdata[447 : 384];
  assign _zz_sram_0_banks_6_bank_port_1 = sram_0_ports_cmd_payload_wstrb[55 : 48];
  assign _zz_sram_0_banks_6_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[6]);
  assign _zz_sram_0_banks_7_bank_port = sram_0_ports_cmd_payload_wdata[511 : 448];
  assign _zz_sram_0_banks_7_bank_port_1 = sram_0_ports_cmd_payload_wstrb[63 : 56];
  assign _zz_sram_0_banks_7_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[7]);
  assign _zz_sram_1_banks_0_bank_port = sram_1_ports_cmd_payload_wdata[63 : 0];
  assign _zz_sram_1_banks_0_bank_port_1 = sram_1_ports_cmd_payload_wstrb[7 : 0];
  assign _zz_sram_1_banks_0_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[0]);
  assign _zz_sram_1_banks_1_bank_port = sram_1_ports_cmd_payload_wdata[127 : 64];
  assign _zz_sram_1_banks_1_bank_port_1 = sram_1_ports_cmd_payload_wstrb[15 : 8];
  assign _zz_sram_1_banks_1_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[1]);
  assign _zz_sram_1_banks_2_bank_port = sram_1_ports_cmd_payload_wdata[191 : 128];
  assign _zz_sram_1_banks_2_bank_port_1 = sram_1_ports_cmd_payload_wstrb[23 : 16];
  assign _zz_sram_1_banks_2_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[2]);
  assign _zz_sram_1_banks_3_bank_port = sram_1_ports_cmd_payload_wdata[255 : 192];
  assign _zz_sram_1_banks_3_bank_port_1 = sram_1_ports_cmd_payload_wstrb[31 : 24];
  assign _zz_sram_1_banks_3_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[3]);
  assign _zz_sram_1_banks_4_bank_port = sram_1_ports_cmd_payload_wdata[319 : 256];
  assign _zz_sram_1_banks_4_bank_port_1 = sram_1_ports_cmd_payload_wstrb[39 : 32];
  assign _zz_sram_1_banks_4_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[4]);
  assign _zz_sram_1_banks_5_bank_port = sram_1_ports_cmd_payload_wdata[383 : 320];
  assign _zz_sram_1_banks_5_bank_port_1 = sram_1_ports_cmd_payload_wstrb[47 : 40];
  assign _zz_sram_1_banks_5_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[5]);
  assign _zz_sram_1_banks_6_bank_port = sram_1_ports_cmd_payload_wdata[447 : 384];
  assign _zz_sram_1_banks_6_bank_port_1 = sram_1_ports_cmd_payload_wstrb[55 : 48];
  assign _zz_sram_1_banks_6_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[6]);
  assign _zz_sram_1_banks_7_bank_port = sram_1_ports_cmd_payload_wdata[511 : 448];
  assign _zz_sram_1_banks_7_bank_port_1 = sram_1_ports_cmd_payload_wstrb[63 : 56];
  assign _zz_sram_1_banks_7_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[7]);
  assign _zz_sram_2_banks_0_bank_port = sram_2_ports_cmd_payload_wdata[63 : 0];
  assign _zz_sram_2_banks_0_bank_port_1 = sram_2_ports_cmd_payload_wstrb[7 : 0];
  assign _zz_sram_2_banks_0_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[0]);
  assign _zz_sram_2_banks_1_bank_port = sram_2_ports_cmd_payload_wdata[127 : 64];
  assign _zz_sram_2_banks_1_bank_port_1 = sram_2_ports_cmd_payload_wstrb[15 : 8];
  assign _zz_sram_2_banks_1_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[1]);
  assign _zz_sram_2_banks_2_bank_port = sram_2_ports_cmd_payload_wdata[191 : 128];
  assign _zz_sram_2_banks_2_bank_port_1 = sram_2_ports_cmd_payload_wstrb[23 : 16];
  assign _zz_sram_2_banks_2_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[2]);
  assign _zz_sram_2_banks_3_bank_port = sram_2_ports_cmd_payload_wdata[255 : 192];
  assign _zz_sram_2_banks_3_bank_port_1 = sram_2_ports_cmd_payload_wstrb[31 : 24];
  assign _zz_sram_2_banks_3_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[3]);
  assign _zz_sram_2_banks_4_bank_port = sram_2_ports_cmd_payload_wdata[319 : 256];
  assign _zz_sram_2_banks_4_bank_port_1 = sram_2_ports_cmd_payload_wstrb[39 : 32];
  assign _zz_sram_2_banks_4_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[4]);
  assign _zz_sram_2_banks_5_bank_port = sram_2_ports_cmd_payload_wdata[383 : 320];
  assign _zz_sram_2_banks_5_bank_port_1 = sram_2_ports_cmd_payload_wstrb[47 : 40];
  assign _zz_sram_2_banks_5_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[5]);
  assign _zz_sram_2_banks_6_bank_port = sram_2_ports_cmd_payload_wdata[447 : 384];
  assign _zz_sram_2_banks_6_bank_port_1 = sram_2_ports_cmd_payload_wstrb[55 : 48];
  assign _zz_sram_2_banks_6_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[6]);
  assign _zz_sram_2_banks_7_bank_port = sram_2_ports_cmd_payload_wdata[511 : 448];
  assign _zz_sram_2_banks_7_bank_port_1 = sram_2_ports_cmd_payload_wstrb[63 : 56];
  assign _zz_sram_2_banks_7_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[7]);
  assign _zz_sram_3_banks_0_bank_port = sram_3_ports_cmd_payload_wdata[63 : 0];
  assign _zz_sram_3_banks_0_bank_port_1 = sram_3_ports_cmd_payload_wstrb[7 : 0];
  assign _zz_sram_3_banks_0_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[0]);
  assign _zz_sram_3_banks_1_bank_port = sram_3_ports_cmd_payload_wdata[127 : 64];
  assign _zz_sram_3_banks_1_bank_port_1 = sram_3_ports_cmd_payload_wstrb[15 : 8];
  assign _zz_sram_3_banks_1_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[1]);
  assign _zz_sram_3_banks_2_bank_port = sram_3_ports_cmd_payload_wdata[191 : 128];
  assign _zz_sram_3_banks_2_bank_port_1 = sram_3_ports_cmd_payload_wstrb[23 : 16];
  assign _zz_sram_3_banks_2_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[2]);
  assign _zz_sram_3_banks_3_bank_port = sram_3_ports_cmd_payload_wdata[255 : 192];
  assign _zz_sram_3_banks_3_bank_port_1 = sram_3_ports_cmd_payload_wstrb[31 : 24];
  assign _zz_sram_3_banks_3_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[3]);
  assign _zz_sram_3_banks_4_bank_port = sram_3_ports_cmd_payload_wdata[319 : 256];
  assign _zz_sram_3_banks_4_bank_port_1 = sram_3_ports_cmd_payload_wstrb[39 : 32];
  assign _zz_sram_3_banks_4_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[4]);
  assign _zz_sram_3_banks_5_bank_port = sram_3_ports_cmd_payload_wdata[383 : 320];
  assign _zz_sram_3_banks_5_bank_port_1 = sram_3_ports_cmd_payload_wstrb[47 : 40];
  assign _zz_sram_3_banks_5_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[5]);
  assign _zz_sram_3_banks_6_bank_port = sram_3_ports_cmd_payload_wdata[447 : 384];
  assign _zz_sram_3_banks_6_bank_port_1 = sram_3_ports_cmd_payload_wstrb[55 : 48];
  assign _zz_sram_3_banks_6_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[6]);
  assign _zz_sram_3_banks_7_bank_port = sram_3_ports_cmd_payload_wdata[511 : 448];
  assign _zz_sram_3_banks_7_bank_port_1 = sram_3_ports_cmd_payload_wstrb[63 : 56];
  assign _zz_sram_3_banks_7_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[7]);
  always @(posedge io_axiClk) begin
    if(_zz_sram_0_banks_0_bank_port_1[0] && _zz_sram_0_banks_0_bank_port_2) begin
      sram_0_banks_0_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_0_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_0_bank_port_1[1] && _zz_sram_0_banks_0_bank_port_2) begin
      sram_0_banks_0_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_0_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_0_bank_port_1[2] && _zz_sram_0_banks_0_bank_port_2) begin
      sram_0_banks_0_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_0_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_0_bank_port_1[3] && _zz_sram_0_banks_0_bank_port_2) begin
      sram_0_banks_0_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_0_bank_port[31 : 24];
    end
    if(_zz_sram_0_banks_0_bank_port_1[4] && _zz_sram_0_banks_0_bank_port_2) begin
      sram_0_banks_0_bank_symbol4[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_0_bank_port[39 : 32];
    end
    if(_zz_sram_0_banks_0_bank_port_1[5] && _zz_sram_0_banks_0_bank_port_2) begin
      sram_0_banks_0_bank_symbol5[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_0_bank_port[47 : 40];
    end
    if(_zz_sram_0_banks_0_bank_port_1[6] && _zz_sram_0_banks_0_bank_port_2) begin
      sram_0_banks_0_bank_symbol6[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_0_bank_port[55 : 48];
    end
    if(_zz_sram_0_banks_0_bank_port_1[7] && _zz_sram_0_banks_0_bank_port_2) begin
      sram_0_banks_0_bank_symbol7[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_0_bank_port[63 : 56];
    end
  end

  assign _zz_sram_0_banks_0_bank_port1[7 : 0] = sram_0_banks_0_bank_symbol0[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_0_bank_port1[15 : 8] = sram_0_banks_0_bank_symbol1[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_0_bank_port1[23 : 16] = sram_0_banks_0_bank_symbol2[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_0_bank_port1[31 : 24] = sram_0_banks_0_bank_symbol3[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_0_bank_port1[39 : 32] = sram_0_banks_0_bank_symbol4[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_0_bank_port1[47 : 40] = sram_0_banks_0_bank_symbol5[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_0_bank_port1[55 : 48] = sram_0_banks_0_bank_symbol6[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_0_bank_port1[63 : 56] = sram_0_banks_0_bank_symbol7[sram_0_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_0_banks_1_bank_port_1[0] && _zz_sram_0_banks_1_bank_port_2) begin
      sram_0_banks_1_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_1_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_1_bank_port_1[1] && _zz_sram_0_banks_1_bank_port_2) begin
      sram_0_banks_1_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_1_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_1_bank_port_1[2] && _zz_sram_0_banks_1_bank_port_2) begin
      sram_0_banks_1_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_1_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_1_bank_port_1[3] && _zz_sram_0_banks_1_bank_port_2) begin
      sram_0_banks_1_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_1_bank_port[31 : 24];
    end
    if(_zz_sram_0_banks_1_bank_port_1[4] && _zz_sram_0_banks_1_bank_port_2) begin
      sram_0_banks_1_bank_symbol4[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_1_bank_port[39 : 32];
    end
    if(_zz_sram_0_banks_1_bank_port_1[5] && _zz_sram_0_banks_1_bank_port_2) begin
      sram_0_banks_1_bank_symbol5[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_1_bank_port[47 : 40];
    end
    if(_zz_sram_0_banks_1_bank_port_1[6] && _zz_sram_0_banks_1_bank_port_2) begin
      sram_0_banks_1_bank_symbol6[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_1_bank_port[55 : 48];
    end
    if(_zz_sram_0_banks_1_bank_port_1[7] && _zz_sram_0_banks_1_bank_port_2) begin
      sram_0_banks_1_bank_symbol7[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_1_bank_port[63 : 56];
    end
  end

  assign _zz_sram_0_banks_1_bank_port1[7 : 0] = sram_0_banks_1_bank_symbol0[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_1_bank_port1[15 : 8] = sram_0_banks_1_bank_symbol1[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_1_bank_port1[23 : 16] = sram_0_banks_1_bank_symbol2[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_1_bank_port1[31 : 24] = sram_0_banks_1_bank_symbol3[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_1_bank_port1[39 : 32] = sram_0_banks_1_bank_symbol4[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_1_bank_port1[47 : 40] = sram_0_banks_1_bank_symbol5[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_1_bank_port1[55 : 48] = sram_0_banks_1_bank_symbol6[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_1_bank_port1[63 : 56] = sram_0_banks_1_bank_symbol7[sram_0_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_0_banks_2_bank_port_1[0] && _zz_sram_0_banks_2_bank_port_2) begin
      sram_0_banks_2_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_2_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_2_bank_port_1[1] && _zz_sram_0_banks_2_bank_port_2) begin
      sram_0_banks_2_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_2_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_2_bank_port_1[2] && _zz_sram_0_banks_2_bank_port_2) begin
      sram_0_banks_2_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_2_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_2_bank_port_1[3] && _zz_sram_0_banks_2_bank_port_2) begin
      sram_0_banks_2_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_2_bank_port[31 : 24];
    end
    if(_zz_sram_0_banks_2_bank_port_1[4] && _zz_sram_0_banks_2_bank_port_2) begin
      sram_0_banks_2_bank_symbol4[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_2_bank_port[39 : 32];
    end
    if(_zz_sram_0_banks_2_bank_port_1[5] && _zz_sram_0_banks_2_bank_port_2) begin
      sram_0_banks_2_bank_symbol5[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_2_bank_port[47 : 40];
    end
    if(_zz_sram_0_banks_2_bank_port_1[6] && _zz_sram_0_banks_2_bank_port_2) begin
      sram_0_banks_2_bank_symbol6[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_2_bank_port[55 : 48];
    end
    if(_zz_sram_0_banks_2_bank_port_1[7] && _zz_sram_0_banks_2_bank_port_2) begin
      sram_0_banks_2_bank_symbol7[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_2_bank_port[63 : 56];
    end
  end

  assign _zz_sram_0_banks_2_bank_port1[7 : 0] = sram_0_banks_2_bank_symbol0[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_2_bank_port1[15 : 8] = sram_0_banks_2_bank_symbol1[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_2_bank_port1[23 : 16] = sram_0_banks_2_bank_symbol2[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_2_bank_port1[31 : 24] = sram_0_banks_2_bank_symbol3[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_2_bank_port1[39 : 32] = sram_0_banks_2_bank_symbol4[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_2_bank_port1[47 : 40] = sram_0_banks_2_bank_symbol5[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_2_bank_port1[55 : 48] = sram_0_banks_2_bank_symbol6[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_2_bank_port1[63 : 56] = sram_0_banks_2_bank_symbol7[sram_0_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_0_banks_3_bank_port_1[0] && _zz_sram_0_banks_3_bank_port_2) begin
      sram_0_banks_3_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_3_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_3_bank_port_1[1] && _zz_sram_0_banks_3_bank_port_2) begin
      sram_0_banks_3_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_3_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_3_bank_port_1[2] && _zz_sram_0_banks_3_bank_port_2) begin
      sram_0_banks_3_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_3_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_3_bank_port_1[3] && _zz_sram_0_banks_3_bank_port_2) begin
      sram_0_banks_3_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_3_bank_port[31 : 24];
    end
    if(_zz_sram_0_banks_3_bank_port_1[4] && _zz_sram_0_banks_3_bank_port_2) begin
      sram_0_banks_3_bank_symbol4[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_3_bank_port[39 : 32];
    end
    if(_zz_sram_0_banks_3_bank_port_1[5] && _zz_sram_0_banks_3_bank_port_2) begin
      sram_0_banks_3_bank_symbol5[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_3_bank_port[47 : 40];
    end
    if(_zz_sram_0_banks_3_bank_port_1[6] && _zz_sram_0_banks_3_bank_port_2) begin
      sram_0_banks_3_bank_symbol6[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_3_bank_port[55 : 48];
    end
    if(_zz_sram_0_banks_3_bank_port_1[7] && _zz_sram_0_banks_3_bank_port_2) begin
      sram_0_banks_3_bank_symbol7[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_3_bank_port[63 : 56];
    end
  end

  assign _zz_sram_0_banks_3_bank_port1[7 : 0] = sram_0_banks_3_bank_symbol0[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_3_bank_port1[15 : 8] = sram_0_banks_3_bank_symbol1[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_3_bank_port1[23 : 16] = sram_0_banks_3_bank_symbol2[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_3_bank_port1[31 : 24] = sram_0_banks_3_bank_symbol3[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_3_bank_port1[39 : 32] = sram_0_banks_3_bank_symbol4[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_3_bank_port1[47 : 40] = sram_0_banks_3_bank_symbol5[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_3_bank_port1[55 : 48] = sram_0_banks_3_bank_symbol6[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_3_bank_port1[63 : 56] = sram_0_banks_3_bank_symbol7[sram_0_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_0_banks_4_bank_port_1[0] && _zz_sram_0_banks_4_bank_port_2) begin
      sram_0_banks_4_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_4_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_4_bank_port_1[1] && _zz_sram_0_banks_4_bank_port_2) begin
      sram_0_banks_4_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_4_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_4_bank_port_1[2] && _zz_sram_0_banks_4_bank_port_2) begin
      sram_0_banks_4_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_4_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_4_bank_port_1[3] && _zz_sram_0_banks_4_bank_port_2) begin
      sram_0_banks_4_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_4_bank_port[31 : 24];
    end
    if(_zz_sram_0_banks_4_bank_port_1[4] && _zz_sram_0_banks_4_bank_port_2) begin
      sram_0_banks_4_bank_symbol4[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_4_bank_port[39 : 32];
    end
    if(_zz_sram_0_banks_4_bank_port_1[5] && _zz_sram_0_banks_4_bank_port_2) begin
      sram_0_banks_4_bank_symbol5[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_4_bank_port[47 : 40];
    end
    if(_zz_sram_0_banks_4_bank_port_1[6] && _zz_sram_0_banks_4_bank_port_2) begin
      sram_0_banks_4_bank_symbol6[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_4_bank_port[55 : 48];
    end
    if(_zz_sram_0_banks_4_bank_port_1[7] && _zz_sram_0_banks_4_bank_port_2) begin
      sram_0_banks_4_bank_symbol7[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_4_bank_port[63 : 56];
    end
  end

  assign _zz_sram_0_banks_4_bank_port1[7 : 0] = sram_0_banks_4_bank_symbol0[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_4_bank_port1[15 : 8] = sram_0_banks_4_bank_symbol1[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_4_bank_port1[23 : 16] = sram_0_banks_4_bank_symbol2[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_4_bank_port1[31 : 24] = sram_0_banks_4_bank_symbol3[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_4_bank_port1[39 : 32] = sram_0_banks_4_bank_symbol4[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_4_bank_port1[47 : 40] = sram_0_banks_4_bank_symbol5[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_4_bank_port1[55 : 48] = sram_0_banks_4_bank_symbol6[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_4_bank_port1[63 : 56] = sram_0_banks_4_bank_symbol7[sram_0_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_0_banks_5_bank_port_1[0] && _zz_sram_0_banks_5_bank_port_2) begin
      sram_0_banks_5_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_5_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_5_bank_port_1[1] && _zz_sram_0_banks_5_bank_port_2) begin
      sram_0_banks_5_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_5_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_5_bank_port_1[2] && _zz_sram_0_banks_5_bank_port_2) begin
      sram_0_banks_5_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_5_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_5_bank_port_1[3] && _zz_sram_0_banks_5_bank_port_2) begin
      sram_0_banks_5_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_5_bank_port[31 : 24];
    end
    if(_zz_sram_0_banks_5_bank_port_1[4] && _zz_sram_0_banks_5_bank_port_2) begin
      sram_0_banks_5_bank_symbol4[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_5_bank_port[39 : 32];
    end
    if(_zz_sram_0_banks_5_bank_port_1[5] && _zz_sram_0_banks_5_bank_port_2) begin
      sram_0_banks_5_bank_symbol5[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_5_bank_port[47 : 40];
    end
    if(_zz_sram_0_banks_5_bank_port_1[6] && _zz_sram_0_banks_5_bank_port_2) begin
      sram_0_banks_5_bank_symbol6[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_5_bank_port[55 : 48];
    end
    if(_zz_sram_0_banks_5_bank_port_1[7] && _zz_sram_0_banks_5_bank_port_2) begin
      sram_0_banks_5_bank_symbol7[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_5_bank_port[63 : 56];
    end
  end

  assign _zz_sram_0_banks_5_bank_port1[7 : 0] = sram_0_banks_5_bank_symbol0[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_5_bank_port1[15 : 8] = sram_0_banks_5_bank_symbol1[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_5_bank_port1[23 : 16] = sram_0_banks_5_bank_symbol2[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_5_bank_port1[31 : 24] = sram_0_banks_5_bank_symbol3[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_5_bank_port1[39 : 32] = sram_0_banks_5_bank_symbol4[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_5_bank_port1[47 : 40] = sram_0_banks_5_bank_symbol5[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_5_bank_port1[55 : 48] = sram_0_banks_5_bank_symbol6[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_5_bank_port1[63 : 56] = sram_0_banks_5_bank_symbol7[sram_0_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_0_banks_6_bank_port_1[0] && _zz_sram_0_banks_6_bank_port_2) begin
      sram_0_banks_6_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_6_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_6_bank_port_1[1] && _zz_sram_0_banks_6_bank_port_2) begin
      sram_0_banks_6_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_6_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_6_bank_port_1[2] && _zz_sram_0_banks_6_bank_port_2) begin
      sram_0_banks_6_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_6_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_6_bank_port_1[3] && _zz_sram_0_banks_6_bank_port_2) begin
      sram_0_banks_6_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_6_bank_port[31 : 24];
    end
    if(_zz_sram_0_banks_6_bank_port_1[4] && _zz_sram_0_banks_6_bank_port_2) begin
      sram_0_banks_6_bank_symbol4[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_6_bank_port[39 : 32];
    end
    if(_zz_sram_0_banks_6_bank_port_1[5] && _zz_sram_0_banks_6_bank_port_2) begin
      sram_0_banks_6_bank_symbol5[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_6_bank_port[47 : 40];
    end
    if(_zz_sram_0_banks_6_bank_port_1[6] && _zz_sram_0_banks_6_bank_port_2) begin
      sram_0_banks_6_bank_symbol6[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_6_bank_port[55 : 48];
    end
    if(_zz_sram_0_banks_6_bank_port_1[7] && _zz_sram_0_banks_6_bank_port_2) begin
      sram_0_banks_6_bank_symbol7[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_6_bank_port[63 : 56];
    end
  end

  assign _zz_sram_0_banks_6_bank_port1[7 : 0] = sram_0_banks_6_bank_symbol0[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_6_bank_port1[15 : 8] = sram_0_banks_6_bank_symbol1[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_6_bank_port1[23 : 16] = sram_0_banks_6_bank_symbol2[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_6_bank_port1[31 : 24] = sram_0_banks_6_bank_symbol3[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_6_bank_port1[39 : 32] = sram_0_banks_6_bank_symbol4[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_6_bank_port1[47 : 40] = sram_0_banks_6_bank_symbol5[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_6_bank_port1[55 : 48] = sram_0_banks_6_bank_symbol6[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_6_bank_port1[63 : 56] = sram_0_banks_6_bank_symbol7[sram_0_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_0_banks_7_bank_port_1[0] && _zz_sram_0_banks_7_bank_port_2) begin
      sram_0_banks_7_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_7_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_7_bank_port_1[1] && _zz_sram_0_banks_7_bank_port_2) begin
      sram_0_banks_7_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_7_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_7_bank_port_1[2] && _zz_sram_0_banks_7_bank_port_2) begin
      sram_0_banks_7_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_7_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_7_bank_port_1[3] && _zz_sram_0_banks_7_bank_port_2) begin
      sram_0_banks_7_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_7_bank_port[31 : 24];
    end
    if(_zz_sram_0_banks_7_bank_port_1[4] && _zz_sram_0_banks_7_bank_port_2) begin
      sram_0_banks_7_bank_symbol4[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_7_bank_port[39 : 32];
    end
    if(_zz_sram_0_banks_7_bank_port_1[5] && _zz_sram_0_banks_7_bank_port_2) begin
      sram_0_banks_7_bank_symbol5[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_7_bank_port[47 : 40];
    end
    if(_zz_sram_0_banks_7_bank_port_1[6] && _zz_sram_0_banks_7_bank_port_2) begin
      sram_0_banks_7_bank_symbol6[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_7_bank_port[55 : 48];
    end
    if(_zz_sram_0_banks_7_bank_port_1[7] && _zz_sram_0_banks_7_bank_port_2) begin
      sram_0_banks_7_bank_symbol7[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_7_bank_port[63 : 56];
    end
  end

  assign _zz_sram_0_banks_7_bank_port1[7 : 0] = sram_0_banks_7_bank_symbol0[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_7_bank_port1[15 : 8] = sram_0_banks_7_bank_symbol1[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_7_bank_port1[23 : 16] = sram_0_banks_7_bank_symbol2[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_7_bank_port1[31 : 24] = sram_0_banks_7_bank_symbol3[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_7_bank_port1[39 : 32] = sram_0_banks_7_bank_symbol4[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_7_bank_port1[47 : 40] = sram_0_banks_7_bank_symbol5[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_7_bank_port1[55 : 48] = sram_0_banks_7_bank_symbol6[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_7_bank_port1[63 : 56] = sram_0_banks_7_bank_symbol7[sram_0_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_1_banks_0_bank_port_1[0] && _zz_sram_1_banks_0_bank_port_2) begin
      sram_1_banks_0_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_0_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_0_bank_port_1[1] && _zz_sram_1_banks_0_bank_port_2) begin
      sram_1_banks_0_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_0_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_0_bank_port_1[2] && _zz_sram_1_banks_0_bank_port_2) begin
      sram_1_banks_0_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_0_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_0_bank_port_1[3] && _zz_sram_1_banks_0_bank_port_2) begin
      sram_1_banks_0_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_0_bank_port[31 : 24];
    end
    if(_zz_sram_1_banks_0_bank_port_1[4] && _zz_sram_1_banks_0_bank_port_2) begin
      sram_1_banks_0_bank_symbol4[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_0_bank_port[39 : 32];
    end
    if(_zz_sram_1_banks_0_bank_port_1[5] && _zz_sram_1_banks_0_bank_port_2) begin
      sram_1_banks_0_bank_symbol5[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_0_bank_port[47 : 40];
    end
    if(_zz_sram_1_banks_0_bank_port_1[6] && _zz_sram_1_banks_0_bank_port_2) begin
      sram_1_banks_0_bank_symbol6[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_0_bank_port[55 : 48];
    end
    if(_zz_sram_1_banks_0_bank_port_1[7] && _zz_sram_1_banks_0_bank_port_2) begin
      sram_1_banks_0_bank_symbol7[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_0_bank_port[63 : 56];
    end
  end

  assign _zz_sram_1_banks_0_bank_port1[7 : 0] = sram_1_banks_0_bank_symbol0[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_0_bank_port1[15 : 8] = sram_1_banks_0_bank_symbol1[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_0_bank_port1[23 : 16] = sram_1_banks_0_bank_symbol2[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_0_bank_port1[31 : 24] = sram_1_banks_0_bank_symbol3[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_0_bank_port1[39 : 32] = sram_1_banks_0_bank_symbol4[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_0_bank_port1[47 : 40] = sram_1_banks_0_bank_symbol5[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_0_bank_port1[55 : 48] = sram_1_banks_0_bank_symbol6[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_0_bank_port1[63 : 56] = sram_1_banks_0_bank_symbol7[sram_1_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_1_banks_1_bank_port_1[0] && _zz_sram_1_banks_1_bank_port_2) begin
      sram_1_banks_1_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_1_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_1_bank_port_1[1] && _zz_sram_1_banks_1_bank_port_2) begin
      sram_1_banks_1_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_1_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_1_bank_port_1[2] && _zz_sram_1_banks_1_bank_port_2) begin
      sram_1_banks_1_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_1_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_1_bank_port_1[3] && _zz_sram_1_banks_1_bank_port_2) begin
      sram_1_banks_1_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_1_bank_port[31 : 24];
    end
    if(_zz_sram_1_banks_1_bank_port_1[4] && _zz_sram_1_banks_1_bank_port_2) begin
      sram_1_banks_1_bank_symbol4[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_1_bank_port[39 : 32];
    end
    if(_zz_sram_1_banks_1_bank_port_1[5] && _zz_sram_1_banks_1_bank_port_2) begin
      sram_1_banks_1_bank_symbol5[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_1_bank_port[47 : 40];
    end
    if(_zz_sram_1_banks_1_bank_port_1[6] && _zz_sram_1_banks_1_bank_port_2) begin
      sram_1_banks_1_bank_symbol6[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_1_bank_port[55 : 48];
    end
    if(_zz_sram_1_banks_1_bank_port_1[7] && _zz_sram_1_banks_1_bank_port_2) begin
      sram_1_banks_1_bank_symbol7[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_1_bank_port[63 : 56];
    end
  end

  assign _zz_sram_1_banks_1_bank_port1[7 : 0] = sram_1_banks_1_bank_symbol0[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_1_bank_port1[15 : 8] = sram_1_banks_1_bank_symbol1[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_1_bank_port1[23 : 16] = sram_1_banks_1_bank_symbol2[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_1_bank_port1[31 : 24] = sram_1_banks_1_bank_symbol3[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_1_bank_port1[39 : 32] = sram_1_banks_1_bank_symbol4[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_1_bank_port1[47 : 40] = sram_1_banks_1_bank_symbol5[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_1_bank_port1[55 : 48] = sram_1_banks_1_bank_symbol6[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_1_bank_port1[63 : 56] = sram_1_banks_1_bank_symbol7[sram_1_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_1_banks_2_bank_port_1[0] && _zz_sram_1_banks_2_bank_port_2) begin
      sram_1_banks_2_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_2_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_2_bank_port_1[1] && _zz_sram_1_banks_2_bank_port_2) begin
      sram_1_banks_2_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_2_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_2_bank_port_1[2] && _zz_sram_1_banks_2_bank_port_2) begin
      sram_1_banks_2_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_2_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_2_bank_port_1[3] && _zz_sram_1_banks_2_bank_port_2) begin
      sram_1_banks_2_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_2_bank_port[31 : 24];
    end
    if(_zz_sram_1_banks_2_bank_port_1[4] && _zz_sram_1_banks_2_bank_port_2) begin
      sram_1_banks_2_bank_symbol4[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_2_bank_port[39 : 32];
    end
    if(_zz_sram_1_banks_2_bank_port_1[5] && _zz_sram_1_banks_2_bank_port_2) begin
      sram_1_banks_2_bank_symbol5[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_2_bank_port[47 : 40];
    end
    if(_zz_sram_1_banks_2_bank_port_1[6] && _zz_sram_1_banks_2_bank_port_2) begin
      sram_1_banks_2_bank_symbol6[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_2_bank_port[55 : 48];
    end
    if(_zz_sram_1_banks_2_bank_port_1[7] && _zz_sram_1_banks_2_bank_port_2) begin
      sram_1_banks_2_bank_symbol7[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_2_bank_port[63 : 56];
    end
  end

  assign _zz_sram_1_banks_2_bank_port1[7 : 0] = sram_1_banks_2_bank_symbol0[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_2_bank_port1[15 : 8] = sram_1_banks_2_bank_symbol1[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_2_bank_port1[23 : 16] = sram_1_banks_2_bank_symbol2[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_2_bank_port1[31 : 24] = sram_1_banks_2_bank_symbol3[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_2_bank_port1[39 : 32] = sram_1_banks_2_bank_symbol4[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_2_bank_port1[47 : 40] = sram_1_banks_2_bank_symbol5[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_2_bank_port1[55 : 48] = sram_1_banks_2_bank_symbol6[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_2_bank_port1[63 : 56] = sram_1_banks_2_bank_symbol7[sram_1_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_1_banks_3_bank_port_1[0] && _zz_sram_1_banks_3_bank_port_2) begin
      sram_1_banks_3_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_3_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_3_bank_port_1[1] && _zz_sram_1_banks_3_bank_port_2) begin
      sram_1_banks_3_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_3_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_3_bank_port_1[2] && _zz_sram_1_banks_3_bank_port_2) begin
      sram_1_banks_3_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_3_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_3_bank_port_1[3] && _zz_sram_1_banks_3_bank_port_2) begin
      sram_1_banks_3_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_3_bank_port[31 : 24];
    end
    if(_zz_sram_1_banks_3_bank_port_1[4] && _zz_sram_1_banks_3_bank_port_2) begin
      sram_1_banks_3_bank_symbol4[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_3_bank_port[39 : 32];
    end
    if(_zz_sram_1_banks_3_bank_port_1[5] && _zz_sram_1_banks_3_bank_port_2) begin
      sram_1_banks_3_bank_symbol5[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_3_bank_port[47 : 40];
    end
    if(_zz_sram_1_banks_3_bank_port_1[6] && _zz_sram_1_banks_3_bank_port_2) begin
      sram_1_banks_3_bank_symbol6[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_3_bank_port[55 : 48];
    end
    if(_zz_sram_1_banks_3_bank_port_1[7] && _zz_sram_1_banks_3_bank_port_2) begin
      sram_1_banks_3_bank_symbol7[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_3_bank_port[63 : 56];
    end
  end

  assign _zz_sram_1_banks_3_bank_port1[7 : 0] = sram_1_banks_3_bank_symbol0[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_3_bank_port1[15 : 8] = sram_1_banks_3_bank_symbol1[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_3_bank_port1[23 : 16] = sram_1_banks_3_bank_symbol2[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_3_bank_port1[31 : 24] = sram_1_banks_3_bank_symbol3[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_3_bank_port1[39 : 32] = sram_1_banks_3_bank_symbol4[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_3_bank_port1[47 : 40] = sram_1_banks_3_bank_symbol5[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_3_bank_port1[55 : 48] = sram_1_banks_3_bank_symbol6[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_3_bank_port1[63 : 56] = sram_1_banks_3_bank_symbol7[sram_1_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_1_banks_4_bank_port_1[0] && _zz_sram_1_banks_4_bank_port_2) begin
      sram_1_banks_4_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_4_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_4_bank_port_1[1] && _zz_sram_1_banks_4_bank_port_2) begin
      sram_1_banks_4_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_4_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_4_bank_port_1[2] && _zz_sram_1_banks_4_bank_port_2) begin
      sram_1_banks_4_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_4_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_4_bank_port_1[3] && _zz_sram_1_banks_4_bank_port_2) begin
      sram_1_banks_4_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_4_bank_port[31 : 24];
    end
    if(_zz_sram_1_banks_4_bank_port_1[4] && _zz_sram_1_banks_4_bank_port_2) begin
      sram_1_banks_4_bank_symbol4[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_4_bank_port[39 : 32];
    end
    if(_zz_sram_1_banks_4_bank_port_1[5] && _zz_sram_1_banks_4_bank_port_2) begin
      sram_1_banks_4_bank_symbol5[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_4_bank_port[47 : 40];
    end
    if(_zz_sram_1_banks_4_bank_port_1[6] && _zz_sram_1_banks_4_bank_port_2) begin
      sram_1_banks_4_bank_symbol6[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_4_bank_port[55 : 48];
    end
    if(_zz_sram_1_banks_4_bank_port_1[7] && _zz_sram_1_banks_4_bank_port_2) begin
      sram_1_banks_4_bank_symbol7[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_4_bank_port[63 : 56];
    end
  end

  assign _zz_sram_1_banks_4_bank_port1[7 : 0] = sram_1_banks_4_bank_symbol0[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_4_bank_port1[15 : 8] = sram_1_banks_4_bank_symbol1[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_4_bank_port1[23 : 16] = sram_1_banks_4_bank_symbol2[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_4_bank_port1[31 : 24] = sram_1_banks_4_bank_symbol3[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_4_bank_port1[39 : 32] = sram_1_banks_4_bank_symbol4[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_4_bank_port1[47 : 40] = sram_1_banks_4_bank_symbol5[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_4_bank_port1[55 : 48] = sram_1_banks_4_bank_symbol6[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_4_bank_port1[63 : 56] = sram_1_banks_4_bank_symbol7[sram_1_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_1_banks_5_bank_port_1[0] && _zz_sram_1_banks_5_bank_port_2) begin
      sram_1_banks_5_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_5_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_5_bank_port_1[1] && _zz_sram_1_banks_5_bank_port_2) begin
      sram_1_banks_5_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_5_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_5_bank_port_1[2] && _zz_sram_1_banks_5_bank_port_2) begin
      sram_1_banks_5_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_5_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_5_bank_port_1[3] && _zz_sram_1_banks_5_bank_port_2) begin
      sram_1_banks_5_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_5_bank_port[31 : 24];
    end
    if(_zz_sram_1_banks_5_bank_port_1[4] && _zz_sram_1_banks_5_bank_port_2) begin
      sram_1_banks_5_bank_symbol4[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_5_bank_port[39 : 32];
    end
    if(_zz_sram_1_banks_5_bank_port_1[5] && _zz_sram_1_banks_5_bank_port_2) begin
      sram_1_banks_5_bank_symbol5[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_5_bank_port[47 : 40];
    end
    if(_zz_sram_1_banks_5_bank_port_1[6] && _zz_sram_1_banks_5_bank_port_2) begin
      sram_1_banks_5_bank_symbol6[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_5_bank_port[55 : 48];
    end
    if(_zz_sram_1_banks_5_bank_port_1[7] && _zz_sram_1_banks_5_bank_port_2) begin
      sram_1_banks_5_bank_symbol7[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_5_bank_port[63 : 56];
    end
  end

  assign _zz_sram_1_banks_5_bank_port1[7 : 0] = sram_1_banks_5_bank_symbol0[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_5_bank_port1[15 : 8] = sram_1_banks_5_bank_symbol1[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_5_bank_port1[23 : 16] = sram_1_banks_5_bank_symbol2[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_5_bank_port1[31 : 24] = sram_1_banks_5_bank_symbol3[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_5_bank_port1[39 : 32] = sram_1_banks_5_bank_symbol4[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_5_bank_port1[47 : 40] = sram_1_banks_5_bank_symbol5[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_5_bank_port1[55 : 48] = sram_1_banks_5_bank_symbol6[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_5_bank_port1[63 : 56] = sram_1_banks_5_bank_symbol7[sram_1_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_1_banks_6_bank_port_1[0] && _zz_sram_1_banks_6_bank_port_2) begin
      sram_1_banks_6_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_6_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_6_bank_port_1[1] && _zz_sram_1_banks_6_bank_port_2) begin
      sram_1_banks_6_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_6_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_6_bank_port_1[2] && _zz_sram_1_banks_6_bank_port_2) begin
      sram_1_banks_6_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_6_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_6_bank_port_1[3] && _zz_sram_1_banks_6_bank_port_2) begin
      sram_1_banks_6_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_6_bank_port[31 : 24];
    end
    if(_zz_sram_1_banks_6_bank_port_1[4] && _zz_sram_1_banks_6_bank_port_2) begin
      sram_1_banks_6_bank_symbol4[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_6_bank_port[39 : 32];
    end
    if(_zz_sram_1_banks_6_bank_port_1[5] && _zz_sram_1_banks_6_bank_port_2) begin
      sram_1_banks_6_bank_symbol5[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_6_bank_port[47 : 40];
    end
    if(_zz_sram_1_banks_6_bank_port_1[6] && _zz_sram_1_banks_6_bank_port_2) begin
      sram_1_banks_6_bank_symbol6[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_6_bank_port[55 : 48];
    end
    if(_zz_sram_1_banks_6_bank_port_1[7] && _zz_sram_1_banks_6_bank_port_2) begin
      sram_1_banks_6_bank_symbol7[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_6_bank_port[63 : 56];
    end
  end

  assign _zz_sram_1_banks_6_bank_port1[7 : 0] = sram_1_banks_6_bank_symbol0[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_6_bank_port1[15 : 8] = sram_1_banks_6_bank_symbol1[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_6_bank_port1[23 : 16] = sram_1_banks_6_bank_symbol2[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_6_bank_port1[31 : 24] = sram_1_banks_6_bank_symbol3[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_6_bank_port1[39 : 32] = sram_1_banks_6_bank_symbol4[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_6_bank_port1[47 : 40] = sram_1_banks_6_bank_symbol5[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_6_bank_port1[55 : 48] = sram_1_banks_6_bank_symbol6[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_6_bank_port1[63 : 56] = sram_1_banks_6_bank_symbol7[sram_1_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_1_banks_7_bank_port_1[0] && _zz_sram_1_banks_7_bank_port_2) begin
      sram_1_banks_7_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_7_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_7_bank_port_1[1] && _zz_sram_1_banks_7_bank_port_2) begin
      sram_1_banks_7_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_7_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_7_bank_port_1[2] && _zz_sram_1_banks_7_bank_port_2) begin
      sram_1_banks_7_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_7_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_7_bank_port_1[3] && _zz_sram_1_banks_7_bank_port_2) begin
      sram_1_banks_7_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_7_bank_port[31 : 24];
    end
    if(_zz_sram_1_banks_7_bank_port_1[4] && _zz_sram_1_banks_7_bank_port_2) begin
      sram_1_banks_7_bank_symbol4[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_7_bank_port[39 : 32];
    end
    if(_zz_sram_1_banks_7_bank_port_1[5] && _zz_sram_1_banks_7_bank_port_2) begin
      sram_1_banks_7_bank_symbol5[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_7_bank_port[47 : 40];
    end
    if(_zz_sram_1_banks_7_bank_port_1[6] && _zz_sram_1_banks_7_bank_port_2) begin
      sram_1_banks_7_bank_symbol6[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_7_bank_port[55 : 48];
    end
    if(_zz_sram_1_banks_7_bank_port_1[7] && _zz_sram_1_banks_7_bank_port_2) begin
      sram_1_banks_7_bank_symbol7[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_7_bank_port[63 : 56];
    end
  end

  assign _zz_sram_1_banks_7_bank_port1[7 : 0] = sram_1_banks_7_bank_symbol0[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_7_bank_port1[15 : 8] = sram_1_banks_7_bank_symbol1[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_7_bank_port1[23 : 16] = sram_1_banks_7_bank_symbol2[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_7_bank_port1[31 : 24] = sram_1_banks_7_bank_symbol3[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_7_bank_port1[39 : 32] = sram_1_banks_7_bank_symbol4[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_7_bank_port1[47 : 40] = sram_1_banks_7_bank_symbol5[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_7_bank_port1[55 : 48] = sram_1_banks_7_bank_symbol6[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_7_bank_port1[63 : 56] = sram_1_banks_7_bank_symbol7[sram_1_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_2_banks_0_bank_port_1[0] && _zz_sram_2_banks_0_bank_port_2) begin
      sram_2_banks_0_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_0_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_0_bank_port_1[1] && _zz_sram_2_banks_0_bank_port_2) begin
      sram_2_banks_0_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_0_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_0_bank_port_1[2] && _zz_sram_2_banks_0_bank_port_2) begin
      sram_2_banks_0_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_0_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_0_bank_port_1[3] && _zz_sram_2_banks_0_bank_port_2) begin
      sram_2_banks_0_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_0_bank_port[31 : 24];
    end
    if(_zz_sram_2_banks_0_bank_port_1[4] && _zz_sram_2_banks_0_bank_port_2) begin
      sram_2_banks_0_bank_symbol4[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_0_bank_port[39 : 32];
    end
    if(_zz_sram_2_banks_0_bank_port_1[5] && _zz_sram_2_banks_0_bank_port_2) begin
      sram_2_banks_0_bank_symbol5[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_0_bank_port[47 : 40];
    end
    if(_zz_sram_2_banks_0_bank_port_1[6] && _zz_sram_2_banks_0_bank_port_2) begin
      sram_2_banks_0_bank_symbol6[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_0_bank_port[55 : 48];
    end
    if(_zz_sram_2_banks_0_bank_port_1[7] && _zz_sram_2_banks_0_bank_port_2) begin
      sram_2_banks_0_bank_symbol7[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_0_bank_port[63 : 56];
    end
  end

  assign _zz_sram_2_banks_0_bank_port1[7 : 0] = sram_2_banks_0_bank_symbol0[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_0_bank_port1[15 : 8] = sram_2_banks_0_bank_symbol1[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_0_bank_port1[23 : 16] = sram_2_banks_0_bank_symbol2[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_0_bank_port1[31 : 24] = sram_2_banks_0_bank_symbol3[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_0_bank_port1[39 : 32] = sram_2_banks_0_bank_symbol4[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_0_bank_port1[47 : 40] = sram_2_banks_0_bank_symbol5[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_0_bank_port1[55 : 48] = sram_2_banks_0_bank_symbol6[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_0_bank_port1[63 : 56] = sram_2_banks_0_bank_symbol7[sram_2_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_2_banks_1_bank_port_1[0] && _zz_sram_2_banks_1_bank_port_2) begin
      sram_2_banks_1_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_1_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_1_bank_port_1[1] && _zz_sram_2_banks_1_bank_port_2) begin
      sram_2_banks_1_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_1_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_1_bank_port_1[2] && _zz_sram_2_banks_1_bank_port_2) begin
      sram_2_banks_1_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_1_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_1_bank_port_1[3] && _zz_sram_2_banks_1_bank_port_2) begin
      sram_2_banks_1_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_1_bank_port[31 : 24];
    end
    if(_zz_sram_2_banks_1_bank_port_1[4] && _zz_sram_2_banks_1_bank_port_2) begin
      sram_2_banks_1_bank_symbol4[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_1_bank_port[39 : 32];
    end
    if(_zz_sram_2_banks_1_bank_port_1[5] && _zz_sram_2_banks_1_bank_port_2) begin
      sram_2_banks_1_bank_symbol5[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_1_bank_port[47 : 40];
    end
    if(_zz_sram_2_banks_1_bank_port_1[6] && _zz_sram_2_banks_1_bank_port_2) begin
      sram_2_banks_1_bank_symbol6[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_1_bank_port[55 : 48];
    end
    if(_zz_sram_2_banks_1_bank_port_1[7] && _zz_sram_2_banks_1_bank_port_2) begin
      sram_2_banks_1_bank_symbol7[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_1_bank_port[63 : 56];
    end
  end

  assign _zz_sram_2_banks_1_bank_port1[7 : 0] = sram_2_banks_1_bank_symbol0[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_1_bank_port1[15 : 8] = sram_2_banks_1_bank_symbol1[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_1_bank_port1[23 : 16] = sram_2_banks_1_bank_symbol2[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_1_bank_port1[31 : 24] = sram_2_banks_1_bank_symbol3[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_1_bank_port1[39 : 32] = sram_2_banks_1_bank_symbol4[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_1_bank_port1[47 : 40] = sram_2_banks_1_bank_symbol5[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_1_bank_port1[55 : 48] = sram_2_banks_1_bank_symbol6[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_1_bank_port1[63 : 56] = sram_2_banks_1_bank_symbol7[sram_2_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_2_banks_2_bank_port_1[0] && _zz_sram_2_banks_2_bank_port_2) begin
      sram_2_banks_2_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_2_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_2_bank_port_1[1] && _zz_sram_2_banks_2_bank_port_2) begin
      sram_2_banks_2_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_2_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_2_bank_port_1[2] && _zz_sram_2_banks_2_bank_port_2) begin
      sram_2_banks_2_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_2_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_2_bank_port_1[3] && _zz_sram_2_banks_2_bank_port_2) begin
      sram_2_banks_2_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_2_bank_port[31 : 24];
    end
    if(_zz_sram_2_banks_2_bank_port_1[4] && _zz_sram_2_banks_2_bank_port_2) begin
      sram_2_banks_2_bank_symbol4[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_2_bank_port[39 : 32];
    end
    if(_zz_sram_2_banks_2_bank_port_1[5] && _zz_sram_2_banks_2_bank_port_2) begin
      sram_2_banks_2_bank_symbol5[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_2_bank_port[47 : 40];
    end
    if(_zz_sram_2_banks_2_bank_port_1[6] && _zz_sram_2_banks_2_bank_port_2) begin
      sram_2_banks_2_bank_symbol6[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_2_bank_port[55 : 48];
    end
    if(_zz_sram_2_banks_2_bank_port_1[7] && _zz_sram_2_banks_2_bank_port_2) begin
      sram_2_banks_2_bank_symbol7[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_2_bank_port[63 : 56];
    end
  end

  assign _zz_sram_2_banks_2_bank_port1[7 : 0] = sram_2_banks_2_bank_symbol0[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_2_bank_port1[15 : 8] = sram_2_banks_2_bank_symbol1[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_2_bank_port1[23 : 16] = sram_2_banks_2_bank_symbol2[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_2_bank_port1[31 : 24] = sram_2_banks_2_bank_symbol3[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_2_bank_port1[39 : 32] = sram_2_banks_2_bank_symbol4[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_2_bank_port1[47 : 40] = sram_2_banks_2_bank_symbol5[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_2_bank_port1[55 : 48] = sram_2_banks_2_bank_symbol6[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_2_bank_port1[63 : 56] = sram_2_banks_2_bank_symbol7[sram_2_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_2_banks_3_bank_port_1[0] && _zz_sram_2_banks_3_bank_port_2) begin
      sram_2_banks_3_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_3_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_3_bank_port_1[1] && _zz_sram_2_banks_3_bank_port_2) begin
      sram_2_banks_3_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_3_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_3_bank_port_1[2] && _zz_sram_2_banks_3_bank_port_2) begin
      sram_2_banks_3_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_3_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_3_bank_port_1[3] && _zz_sram_2_banks_3_bank_port_2) begin
      sram_2_banks_3_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_3_bank_port[31 : 24];
    end
    if(_zz_sram_2_banks_3_bank_port_1[4] && _zz_sram_2_banks_3_bank_port_2) begin
      sram_2_banks_3_bank_symbol4[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_3_bank_port[39 : 32];
    end
    if(_zz_sram_2_banks_3_bank_port_1[5] && _zz_sram_2_banks_3_bank_port_2) begin
      sram_2_banks_3_bank_symbol5[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_3_bank_port[47 : 40];
    end
    if(_zz_sram_2_banks_3_bank_port_1[6] && _zz_sram_2_banks_3_bank_port_2) begin
      sram_2_banks_3_bank_symbol6[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_3_bank_port[55 : 48];
    end
    if(_zz_sram_2_banks_3_bank_port_1[7] && _zz_sram_2_banks_3_bank_port_2) begin
      sram_2_banks_3_bank_symbol7[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_3_bank_port[63 : 56];
    end
  end

  assign _zz_sram_2_banks_3_bank_port1[7 : 0] = sram_2_banks_3_bank_symbol0[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_3_bank_port1[15 : 8] = sram_2_banks_3_bank_symbol1[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_3_bank_port1[23 : 16] = sram_2_banks_3_bank_symbol2[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_3_bank_port1[31 : 24] = sram_2_banks_3_bank_symbol3[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_3_bank_port1[39 : 32] = sram_2_banks_3_bank_symbol4[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_3_bank_port1[47 : 40] = sram_2_banks_3_bank_symbol5[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_3_bank_port1[55 : 48] = sram_2_banks_3_bank_symbol6[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_3_bank_port1[63 : 56] = sram_2_banks_3_bank_symbol7[sram_2_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_2_banks_4_bank_port_1[0] && _zz_sram_2_banks_4_bank_port_2) begin
      sram_2_banks_4_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_4_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_4_bank_port_1[1] && _zz_sram_2_banks_4_bank_port_2) begin
      sram_2_banks_4_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_4_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_4_bank_port_1[2] && _zz_sram_2_banks_4_bank_port_2) begin
      sram_2_banks_4_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_4_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_4_bank_port_1[3] && _zz_sram_2_banks_4_bank_port_2) begin
      sram_2_banks_4_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_4_bank_port[31 : 24];
    end
    if(_zz_sram_2_banks_4_bank_port_1[4] && _zz_sram_2_banks_4_bank_port_2) begin
      sram_2_banks_4_bank_symbol4[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_4_bank_port[39 : 32];
    end
    if(_zz_sram_2_banks_4_bank_port_1[5] && _zz_sram_2_banks_4_bank_port_2) begin
      sram_2_banks_4_bank_symbol5[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_4_bank_port[47 : 40];
    end
    if(_zz_sram_2_banks_4_bank_port_1[6] && _zz_sram_2_banks_4_bank_port_2) begin
      sram_2_banks_4_bank_symbol6[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_4_bank_port[55 : 48];
    end
    if(_zz_sram_2_banks_4_bank_port_1[7] && _zz_sram_2_banks_4_bank_port_2) begin
      sram_2_banks_4_bank_symbol7[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_4_bank_port[63 : 56];
    end
  end

  assign _zz_sram_2_banks_4_bank_port1[7 : 0] = sram_2_banks_4_bank_symbol0[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_4_bank_port1[15 : 8] = sram_2_banks_4_bank_symbol1[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_4_bank_port1[23 : 16] = sram_2_banks_4_bank_symbol2[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_4_bank_port1[31 : 24] = sram_2_banks_4_bank_symbol3[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_4_bank_port1[39 : 32] = sram_2_banks_4_bank_symbol4[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_4_bank_port1[47 : 40] = sram_2_banks_4_bank_symbol5[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_4_bank_port1[55 : 48] = sram_2_banks_4_bank_symbol6[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_4_bank_port1[63 : 56] = sram_2_banks_4_bank_symbol7[sram_2_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_2_banks_5_bank_port_1[0] && _zz_sram_2_banks_5_bank_port_2) begin
      sram_2_banks_5_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_5_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_5_bank_port_1[1] && _zz_sram_2_banks_5_bank_port_2) begin
      sram_2_banks_5_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_5_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_5_bank_port_1[2] && _zz_sram_2_banks_5_bank_port_2) begin
      sram_2_banks_5_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_5_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_5_bank_port_1[3] && _zz_sram_2_banks_5_bank_port_2) begin
      sram_2_banks_5_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_5_bank_port[31 : 24];
    end
    if(_zz_sram_2_banks_5_bank_port_1[4] && _zz_sram_2_banks_5_bank_port_2) begin
      sram_2_banks_5_bank_symbol4[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_5_bank_port[39 : 32];
    end
    if(_zz_sram_2_banks_5_bank_port_1[5] && _zz_sram_2_banks_5_bank_port_2) begin
      sram_2_banks_5_bank_symbol5[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_5_bank_port[47 : 40];
    end
    if(_zz_sram_2_banks_5_bank_port_1[6] && _zz_sram_2_banks_5_bank_port_2) begin
      sram_2_banks_5_bank_symbol6[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_5_bank_port[55 : 48];
    end
    if(_zz_sram_2_banks_5_bank_port_1[7] && _zz_sram_2_banks_5_bank_port_2) begin
      sram_2_banks_5_bank_symbol7[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_5_bank_port[63 : 56];
    end
  end

  assign _zz_sram_2_banks_5_bank_port1[7 : 0] = sram_2_banks_5_bank_symbol0[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_5_bank_port1[15 : 8] = sram_2_banks_5_bank_symbol1[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_5_bank_port1[23 : 16] = sram_2_banks_5_bank_symbol2[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_5_bank_port1[31 : 24] = sram_2_banks_5_bank_symbol3[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_5_bank_port1[39 : 32] = sram_2_banks_5_bank_symbol4[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_5_bank_port1[47 : 40] = sram_2_banks_5_bank_symbol5[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_5_bank_port1[55 : 48] = sram_2_banks_5_bank_symbol6[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_5_bank_port1[63 : 56] = sram_2_banks_5_bank_symbol7[sram_2_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_2_banks_6_bank_port_1[0] && _zz_sram_2_banks_6_bank_port_2) begin
      sram_2_banks_6_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_6_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_6_bank_port_1[1] && _zz_sram_2_banks_6_bank_port_2) begin
      sram_2_banks_6_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_6_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_6_bank_port_1[2] && _zz_sram_2_banks_6_bank_port_2) begin
      sram_2_banks_6_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_6_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_6_bank_port_1[3] && _zz_sram_2_banks_6_bank_port_2) begin
      sram_2_banks_6_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_6_bank_port[31 : 24];
    end
    if(_zz_sram_2_banks_6_bank_port_1[4] && _zz_sram_2_banks_6_bank_port_2) begin
      sram_2_banks_6_bank_symbol4[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_6_bank_port[39 : 32];
    end
    if(_zz_sram_2_banks_6_bank_port_1[5] && _zz_sram_2_banks_6_bank_port_2) begin
      sram_2_banks_6_bank_symbol5[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_6_bank_port[47 : 40];
    end
    if(_zz_sram_2_banks_6_bank_port_1[6] && _zz_sram_2_banks_6_bank_port_2) begin
      sram_2_banks_6_bank_symbol6[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_6_bank_port[55 : 48];
    end
    if(_zz_sram_2_banks_6_bank_port_1[7] && _zz_sram_2_banks_6_bank_port_2) begin
      sram_2_banks_6_bank_symbol7[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_6_bank_port[63 : 56];
    end
  end

  assign _zz_sram_2_banks_6_bank_port1[7 : 0] = sram_2_banks_6_bank_symbol0[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_6_bank_port1[15 : 8] = sram_2_banks_6_bank_symbol1[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_6_bank_port1[23 : 16] = sram_2_banks_6_bank_symbol2[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_6_bank_port1[31 : 24] = sram_2_banks_6_bank_symbol3[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_6_bank_port1[39 : 32] = sram_2_banks_6_bank_symbol4[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_6_bank_port1[47 : 40] = sram_2_banks_6_bank_symbol5[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_6_bank_port1[55 : 48] = sram_2_banks_6_bank_symbol6[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_6_bank_port1[63 : 56] = sram_2_banks_6_bank_symbol7[sram_2_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_2_banks_7_bank_port_1[0] && _zz_sram_2_banks_7_bank_port_2) begin
      sram_2_banks_7_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_7_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_7_bank_port_1[1] && _zz_sram_2_banks_7_bank_port_2) begin
      sram_2_banks_7_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_7_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_7_bank_port_1[2] && _zz_sram_2_banks_7_bank_port_2) begin
      sram_2_banks_7_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_7_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_7_bank_port_1[3] && _zz_sram_2_banks_7_bank_port_2) begin
      sram_2_banks_7_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_7_bank_port[31 : 24];
    end
    if(_zz_sram_2_banks_7_bank_port_1[4] && _zz_sram_2_banks_7_bank_port_2) begin
      sram_2_banks_7_bank_symbol4[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_7_bank_port[39 : 32];
    end
    if(_zz_sram_2_banks_7_bank_port_1[5] && _zz_sram_2_banks_7_bank_port_2) begin
      sram_2_banks_7_bank_symbol5[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_7_bank_port[47 : 40];
    end
    if(_zz_sram_2_banks_7_bank_port_1[6] && _zz_sram_2_banks_7_bank_port_2) begin
      sram_2_banks_7_bank_symbol6[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_7_bank_port[55 : 48];
    end
    if(_zz_sram_2_banks_7_bank_port_1[7] && _zz_sram_2_banks_7_bank_port_2) begin
      sram_2_banks_7_bank_symbol7[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_7_bank_port[63 : 56];
    end
  end

  assign _zz_sram_2_banks_7_bank_port1[7 : 0] = sram_2_banks_7_bank_symbol0[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_7_bank_port1[15 : 8] = sram_2_banks_7_bank_symbol1[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_7_bank_port1[23 : 16] = sram_2_banks_7_bank_symbol2[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_7_bank_port1[31 : 24] = sram_2_banks_7_bank_symbol3[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_7_bank_port1[39 : 32] = sram_2_banks_7_bank_symbol4[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_7_bank_port1[47 : 40] = sram_2_banks_7_bank_symbol5[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_7_bank_port1[55 : 48] = sram_2_banks_7_bank_symbol6[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_7_bank_port1[63 : 56] = sram_2_banks_7_bank_symbol7[sram_2_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_3_banks_0_bank_port_1[0] && _zz_sram_3_banks_0_bank_port_2) begin
      sram_3_banks_0_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_0_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_0_bank_port_1[1] && _zz_sram_3_banks_0_bank_port_2) begin
      sram_3_banks_0_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_0_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_0_bank_port_1[2] && _zz_sram_3_banks_0_bank_port_2) begin
      sram_3_banks_0_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_0_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_0_bank_port_1[3] && _zz_sram_3_banks_0_bank_port_2) begin
      sram_3_banks_0_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_0_bank_port[31 : 24];
    end
    if(_zz_sram_3_banks_0_bank_port_1[4] && _zz_sram_3_banks_0_bank_port_2) begin
      sram_3_banks_0_bank_symbol4[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_0_bank_port[39 : 32];
    end
    if(_zz_sram_3_banks_0_bank_port_1[5] && _zz_sram_3_banks_0_bank_port_2) begin
      sram_3_banks_0_bank_symbol5[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_0_bank_port[47 : 40];
    end
    if(_zz_sram_3_banks_0_bank_port_1[6] && _zz_sram_3_banks_0_bank_port_2) begin
      sram_3_banks_0_bank_symbol6[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_0_bank_port[55 : 48];
    end
    if(_zz_sram_3_banks_0_bank_port_1[7] && _zz_sram_3_banks_0_bank_port_2) begin
      sram_3_banks_0_bank_symbol7[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_0_bank_port[63 : 56];
    end
  end

  assign _zz_sram_3_banks_0_bank_port1[7 : 0] = sram_3_banks_0_bank_symbol0[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_0_bank_port1[15 : 8] = sram_3_banks_0_bank_symbol1[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_0_bank_port1[23 : 16] = sram_3_banks_0_bank_symbol2[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_0_bank_port1[31 : 24] = sram_3_banks_0_bank_symbol3[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_0_bank_port1[39 : 32] = sram_3_banks_0_bank_symbol4[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_0_bank_port1[47 : 40] = sram_3_banks_0_bank_symbol5[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_0_bank_port1[55 : 48] = sram_3_banks_0_bank_symbol6[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_0_bank_port1[63 : 56] = sram_3_banks_0_bank_symbol7[sram_3_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_3_banks_1_bank_port_1[0] && _zz_sram_3_banks_1_bank_port_2) begin
      sram_3_banks_1_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_1_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_1_bank_port_1[1] && _zz_sram_3_banks_1_bank_port_2) begin
      sram_3_banks_1_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_1_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_1_bank_port_1[2] && _zz_sram_3_banks_1_bank_port_2) begin
      sram_3_banks_1_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_1_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_1_bank_port_1[3] && _zz_sram_3_banks_1_bank_port_2) begin
      sram_3_banks_1_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_1_bank_port[31 : 24];
    end
    if(_zz_sram_3_banks_1_bank_port_1[4] && _zz_sram_3_banks_1_bank_port_2) begin
      sram_3_banks_1_bank_symbol4[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_1_bank_port[39 : 32];
    end
    if(_zz_sram_3_banks_1_bank_port_1[5] && _zz_sram_3_banks_1_bank_port_2) begin
      sram_3_banks_1_bank_symbol5[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_1_bank_port[47 : 40];
    end
    if(_zz_sram_3_banks_1_bank_port_1[6] && _zz_sram_3_banks_1_bank_port_2) begin
      sram_3_banks_1_bank_symbol6[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_1_bank_port[55 : 48];
    end
    if(_zz_sram_3_banks_1_bank_port_1[7] && _zz_sram_3_banks_1_bank_port_2) begin
      sram_3_banks_1_bank_symbol7[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_1_bank_port[63 : 56];
    end
  end

  assign _zz_sram_3_banks_1_bank_port1[7 : 0] = sram_3_banks_1_bank_symbol0[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_1_bank_port1[15 : 8] = sram_3_banks_1_bank_symbol1[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_1_bank_port1[23 : 16] = sram_3_banks_1_bank_symbol2[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_1_bank_port1[31 : 24] = sram_3_banks_1_bank_symbol3[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_1_bank_port1[39 : 32] = sram_3_banks_1_bank_symbol4[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_1_bank_port1[47 : 40] = sram_3_banks_1_bank_symbol5[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_1_bank_port1[55 : 48] = sram_3_banks_1_bank_symbol6[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_1_bank_port1[63 : 56] = sram_3_banks_1_bank_symbol7[sram_3_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_3_banks_2_bank_port_1[0] && _zz_sram_3_banks_2_bank_port_2) begin
      sram_3_banks_2_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_2_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_2_bank_port_1[1] && _zz_sram_3_banks_2_bank_port_2) begin
      sram_3_banks_2_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_2_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_2_bank_port_1[2] && _zz_sram_3_banks_2_bank_port_2) begin
      sram_3_banks_2_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_2_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_2_bank_port_1[3] && _zz_sram_3_banks_2_bank_port_2) begin
      sram_3_banks_2_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_2_bank_port[31 : 24];
    end
    if(_zz_sram_3_banks_2_bank_port_1[4] && _zz_sram_3_banks_2_bank_port_2) begin
      sram_3_banks_2_bank_symbol4[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_2_bank_port[39 : 32];
    end
    if(_zz_sram_3_banks_2_bank_port_1[5] && _zz_sram_3_banks_2_bank_port_2) begin
      sram_3_banks_2_bank_symbol5[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_2_bank_port[47 : 40];
    end
    if(_zz_sram_3_banks_2_bank_port_1[6] && _zz_sram_3_banks_2_bank_port_2) begin
      sram_3_banks_2_bank_symbol6[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_2_bank_port[55 : 48];
    end
    if(_zz_sram_3_banks_2_bank_port_1[7] && _zz_sram_3_banks_2_bank_port_2) begin
      sram_3_banks_2_bank_symbol7[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_2_bank_port[63 : 56];
    end
  end

  assign _zz_sram_3_banks_2_bank_port1[7 : 0] = sram_3_banks_2_bank_symbol0[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_2_bank_port1[15 : 8] = sram_3_banks_2_bank_symbol1[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_2_bank_port1[23 : 16] = sram_3_banks_2_bank_symbol2[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_2_bank_port1[31 : 24] = sram_3_banks_2_bank_symbol3[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_2_bank_port1[39 : 32] = sram_3_banks_2_bank_symbol4[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_2_bank_port1[47 : 40] = sram_3_banks_2_bank_symbol5[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_2_bank_port1[55 : 48] = sram_3_banks_2_bank_symbol6[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_2_bank_port1[63 : 56] = sram_3_banks_2_bank_symbol7[sram_3_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_3_banks_3_bank_port_1[0] && _zz_sram_3_banks_3_bank_port_2) begin
      sram_3_banks_3_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_3_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_3_bank_port_1[1] && _zz_sram_3_banks_3_bank_port_2) begin
      sram_3_banks_3_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_3_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_3_bank_port_1[2] && _zz_sram_3_banks_3_bank_port_2) begin
      sram_3_banks_3_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_3_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_3_bank_port_1[3] && _zz_sram_3_banks_3_bank_port_2) begin
      sram_3_banks_3_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_3_bank_port[31 : 24];
    end
    if(_zz_sram_3_banks_3_bank_port_1[4] && _zz_sram_3_banks_3_bank_port_2) begin
      sram_3_banks_3_bank_symbol4[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_3_bank_port[39 : 32];
    end
    if(_zz_sram_3_banks_3_bank_port_1[5] && _zz_sram_3_banks_3_bank_port_2) begin
      sram_3_banks_3_bank_symbol5[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_3_bank_port[47 : 40];
    end
    if(_zz_sram_3_banks_3_bank_port_1[6] && _zz_sram_3_banks_3_bank_port_2) begin
      sram_3_banks_3_bank_symbol6[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_3_bank_port[55 : 48];
    end
    if(_zz_sram_3_banks_3_bank_port_1[7] && _zz_sram_3_banks_3_bank_port_2) begin
      sram_3_banks_3_bank_symbol7[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_3_bank_port[63 : 56];
    end
  end

  assign _zz_sram_3_banks_3_bank_port1[7 : 0] = sram_3_banks_3_bank_symbol0[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_3_bank_port1[15 : 8] = sram_3_banks_3_bank_symbol1[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_3_bank_port1[23 : 16] = sram_3_banks_3_bank_symbol2[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_3_bank_port1[31 : 24] = sram_3_banks_3_bank_symbol3[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_3_bank_port1[39 : 32] = sram_3_banks_3_bank_symbol4[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_3_bank_port1[47 : 40] = sram_3_banks_3_bank_symbol5[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_3_bank_port1[55 : 48] = sram_3_banks_3_bank_symbol6[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_3_bank_port1[63 : 56] = sram_3_banks_3_bank_symbol7[sram_3_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_3_banks_4_bank_port_1[0] && _zz_sram_3_banks_4_bank_port_2) begin
      sram_3_banks_4_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_4_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_4_bank_port_1[1] && _zz_sram_3_banks_4_bank_port_2) begin
      sram_3_banks_4_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_4_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_4_bank_port_1[2] && _zz_sram_3_banks_4_bank_port_2) begin
      sram_3_banks_4_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_4_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_4_bank_port_1[3] && _zz_sram_3_banks_4_bank_port_2) begin
      sram_3_banks_4_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_4_bank_port[31 : 24];
    end
    if(_zz_sram_3_banks_4_bank_port_1[4] && _zz_sram_3_banks_4_bank_port_2) begin
      sram_3_banks_4_bank_symbol4[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_4_bank_port[39 : 32];
    end
    if(_zz_sram_3_banks_4_bank_port_1[5] && _zz_sram_3_banks_4_bank_port_2) begin
      sram_3_banks_4_bank_symbol5[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_4_bank_port[47 : 40];
    end
    if(_zz_sram_3_banks_4_bank_port_1[6] && _zz_sram_3_banks_4_bank_port_2) begin
      sram_3_banks_4_bank_symbol6[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_4_bank_port[55 : 48];
    end
    if(_zz_sram_3_banks_4_bank_port_1[7] && _zz_sram_3_banks_4_bank_port_2) begin
      sram_3_banks_4_bank_symbol7[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_4_bank_port[63 : 56];
    end
  end

  assign _zz_sram_3_banks_4_bank_port1[7 : 0] = sram_3_banks_4_bank_symbol0[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_4_bank_port1[15 : 8] = sram_3_banks_4_bank_symbol1[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_4_bank_port1[23 : 16] = sram_3_banks_4_bank_symbol2[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_4_bank_port1[31 : 24] = sram_3_banks_4_bank_symbol3[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_4_bank_port1[39 : 32] = sram_3_banks_4_bank_symbol4[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_4_bank_port1[47 : 40] = sram_3_banks_4_bank_symbol5[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_4_bank_port1[55 : 48] = sram_3_banks_4_bank_symbol6[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_4_bank_port1[63 : 56] = sram_3_banks_4_bank_symbol7[sram_3_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_3_banks_5_bank_port_1[0] && _zz_sram_3_banks_5_bank_port_2) begin
      sram_3_banks_5_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_5_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_5_bank_port_1[1] && _zz_sram_3_banks_5_bank_port_2) begin
      sram_3_banks_5_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_5_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_5_bank_port_1[2] && _zz_sram_3_banks_5_bank_port_2) begin
      sram_3_banks_5_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_5_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_5_bank_port_1[3] && _zz_sram_3_banks_5_bank_port_2) begin
      sram_3_banks_5_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_5_bank_port[31 : 24];
    end
    if(_zz_sram_3_banks_5_bank_port_1[4] && _zz_sram_3_banks_5_bank_port_2) begin
      sram_3_banks_5_bank_symbol4[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_5_bank_port[39 : 32];
    end
    if(_zz_sram_3_banks_5_bank_port_1[5] && _zz_sram_3_banks_5_bank_port_2) begin
      sram_3_banks_5_bank_symbol5[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_5_bank_port[47 : 40];
    end
    if(_zz_sram_3_banks_5_bank_port_1[6] && _zz_sram_3_banks_5_bank_port_2) begin
      sram_3_banks_5_bank_symbol6[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_5_bank_port[55 : 48];
    end
    if(_zz_sram_3_banks_5_bank_port_1[7] && _zz_sram_3_banks_5_bank_port_2) begin
      sram_3_banks_5_bank_symbol7[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_5_bank_port[63 : 56];
    end
  end

  assign _zz_sram_3_banks_5_bank_port1[7 : 0] = sram_3_banks_5_bank_symbol0[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_5_bank_port1[15 : 8] = sram_3_banks_5_bank_symbol1[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_5_bank_port1[23 : 16] = sram_3_banks_5_bank_symbol2[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_5_bank_port1[31 : 24] = sram_3_banks_5_bank_symbol3[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_5_bank_port1[39 : 32] = sram_3_banks_5_bank_symbol4[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_5_bank_port1[47 : 40] = sram_3_banks_5_bank_symbol5[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_5_bank_port1[55 : 48] = sram_3_banks_5_bank_symbol6[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_5_bank_port1[63 : 56] = sram_3_banks_5_bank_symbol7[sram_3_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_3_banks_6_bank_port_1[0] && _zz_sram_3_banks_6_bank_port_2) begin
      sram_3_banks_6_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_6_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_6_bank_port_1[1] && _zz_sram_3_banks_6_bank_port_2) begin
      sram_3_banks_6_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_6_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_6_bank_port_1[2] && _zz_sram_3_banks_6_bank_port_2) begin
      sram_3_banks_6_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_6_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_6_bank_port_1[3] && _zz_sram_3_banks_6_bank_port_2) begin
      sram_3_banks_6_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_6_bank_port[31 : 24];
    end
    if(_zz_sram_3_banks_6_bank_port_1[4] && _zz_sram_3_banks_6_bank_port_2) begin
      sram_3_banks_6_bank_symbol4[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_6_bank_port[39 : 32];
    end
    if(_zz_sram_3_banks_6_bank_port_1[5] && _zz_sram_3_banks_6_bank_port_2) begin
      sram_3_banks_6_bank_symbol5[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_6_bank_port[47 : 40];
    end
    if(_zz_sram_3_banks_6_bank_port_1[6] && _zz_sram_3_banks_6_bank_port_2) begin
      sram_3_banks_6_bank_symbol6[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_6_bank_port[55 : 48];
    end
    if(_zz_sram_3_banks_6_bank_port_1[7] && _zz_sram_3_banks_6_bank_port_2) begin
      sram_3_banks_6_bank_symbol7[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_6_bank_port[63 : 56];
    end
  end

  assign _zz_sram_3_banks_6_bank_port1[7 : 0] = sram_3_banks_6_bank_symbol0[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_6_bank_port1[15 : 8] = sram_3_banks_6_bank_symbol1[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_6_bank_port1[23 : 16] = sram_3_banks_6_bank_symbol2[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_6_bank_port1[31 : 24] = sram_3_banks_6_bank_symbol3[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_6_bank_port1[39 : 32] = sram_3_banks_6_bank_symbol4[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_6_bank_port1[47 : 40] = sram_3_banks_6_bank_symbol5[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_6_bank_port1[55 : 48] = sram_3_banks_6_bank_symbol6[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_6_bank_port1[63 : 56] = sram_3_banks_6_bank_symbol7[sram_3_ports_cmd_payload_addr];
  always @(posedge io_axiClk) begin
    if(_zz_sram_3_banks_7_bank_port_1[0] && _zz_sram_3_banks_7_bank_port_2) begin
      sram_3_banks_7_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_7_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_7_bank_port_1[1] && _zz_sram_3_banks_7_bank_port_2) begin
      sram_3_banks_7_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_7_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_7_bank_port_1[2] && _zz_sram_3_banks_7_bank_port_2) begin
      sram_3_banks_7_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_7_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_7_bank_port_1[3] && _zz_sram_3_banks_7_bank_port_2) begin
      sram_3_banks_7_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_7_bank_port[31 : 24];
    end
    if(_zz_sram_3_banks_7_bank_port_1[4] && _zz_sram_3_banks_7_bank_port_2) begin
      sram_3_banks_7_bank_symbol4[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_7_bank_port[39 : 32];
    end
    if(_zz_sram_3_banks_7_bank_port_1[5] && _zz_sram_3_banks_7_bank_port_2) begin
      sram_3_banks_7_bank_symbol5[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_7_bank_port[47 : 40];
    end
    if(_zz_sram_3_banks_7_bank_port_1[6] && _zz_sram_3_banks_7_bank_port_2) begin
      sram_3_banks_7_bank_symbol6[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_7_bank_port[55 : 48];
    end
    if(_zz_sram_3_banks_7_bank_port_1[7] && _zz_sram_3_banks_7_bank_port_2) begin
      sram_3_banks_7_bank_symbol7[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_7_bank_port[63 : 56];
    end
  end

  assign _zz_sram_3_banks_7_bank_port1[7 : 0] = sram_3_banks_7_bank_symbol0[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_7_bank_port1[15 : 8] = sram_3_banks_7_bank_symbol1[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_7_bank_port1[23 : 16] = sram_3_banks_7_bank_symbol2[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_7_bank_port1[31 : 24] = sram_3_banks_7_bank_symbol3[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_7_bank_port1[39 : 32] = sram_3_banks_7_bank_symbol4[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_7_bank_port1[47 : 40] = sram_3_banks_7_bank_symbol5[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_7_bank_port1[55 : 48] = sram_3_banks_7_bank_symbol6[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_7_bank_port1[63 : 56] = sram_3_banks_7_bank_symbol7[sram_3_ports_cmd_payload_addr];
  always @(*) begin
    sram_0_ports_rsp_payload_data[63 : 0] = _zz_sram_0_banks_0_bank_port1;
    sram_0_ports_rsp_payload_data[127 : 64] = _zz_sram_0_banks_1_bank_port1;
    sram_0_ports_rsp_payload_data[191 : 128] = _zz_sram_0_banks_2_bank_port1;
    sram_0_ports_rsp_payload_data[255 : 192] = _zz_sram_0_banks_3_bank_port1;
    sram_0_ports_rsp_payload_data[319 : 256] = _zz_sram_0_banks_4_bank_port1;
    sram_0_ports_rsp_payload_data[383 : 320] = _zz_sram_0_banks_5_bank_port1;
    sram_0_ports_rsp_payload_data[447 : 384] = _zz_sram_0_banks_6_bank_port1;
    sram_0_ports_rsp_payload_data[511 : 448] = _zz_sram_0_banks_7_bank_port1;
  end

  assign when_SramBanks_l75 = (sram_0_ports_cmd_valid && (sram_0_ports_cmd_payload_wen == 8'h0));
  always @(*) begin
    if(when_SramBanks_l75) begin
      _zz_sram_0_ports_rsp_valid = 1'b1;
    end else begin
      _zz_sram_0_ports_rsp_valid = 1'b0;
    end
  end

  assign sram_0_ports_rsp_valid = _zz_sram_0_ports_rsp_valid;
  always @(*) begin
    sram_1_ports_rsp_payload_data[63 : 0] = _zz_sram_1_banks_0_bank_port1;
    sram_1_ports_rsp_payload_data[127 : 64] = _zz_sram_1_banks_1_bank_port1;
    sram_1_ports_rsp_payload_data[191 : 128] = _zz_sram_1_banks_2_bank_port1;
    sram_1_ports_rsp_payload_data[255 : 192] = _zz_sram_1_banks_3_bank_port1;
    sram_1_ports_rsp_payload_data[319 : 256] = _zz_sram_1_banks_4_bank_port1;
    sram_1_ports_rsp_payload_data[383 : 320] = _zz_sram_1_banks_5_bank_port1;
    sram_1_ports_rsp_payload_data[447 : 384] = _zz_sram_1_banks_6_bank_port1;
    sram_1_ports_rsp_payload_data[511 : 448] = _zz_sram_1_banks_7_bank_port1;
  end

  assign when_SramBanks_l75_1 = (sram_1_ports_cmd_valid && (sram_1_ports_cmd_payload_wen == 8'h0));
  always @(*) begin
    if(when_SramBanks_l75_1) begin
      _zz_sram_1_ports_rsp_valid = 1'b1;
    end else begin
      _zz_sram_1_ports_rsp_valid = 1'b0;
    end
  end

  assign sram_1_ports_rsp_valid = _zz_sram_1_ports_rsp_valid;
  always @(*) begin
    sram_2_ports_rsp_payload_data[63 : 0] = _zz_sram_2_banks_0_bank_port1;
    sram_2_ports_rsp_payload_data[127 : 64] = _zz_sram_2_banks_1_bank_port1;
    sram_2_ports_rsp_payload_data[191 : 128] = _zz_sram_2_banks_2_bank_port1;
    sram_2_ports_rsp_payload_data[255 : 192] = _zz_sram_2_banks_3_bank_port1;
    sram_2_ports_rsp_payload_data[319 : 256] = _zz_sram_2_banks_4_bank_port1;
    sram_2_ports_rsp_payload_data[383 : 320] = _zz_sram_2_banks_5_bank_port1;
    sram_2_ports_rsp_payload_data[447 : 384] = _zz_sram_2_banks_6_bank_port1;
    sram_2_ports_rsp_payload_data[511 : 448] = _zz_sram_2_banks_7_bank_port1;
  end

  assign when_SramBanks_l75_2 = (sram_2_ports_cmd_valid && (sram_2_ports_cmd_payload_wen == 8'h0));
  always @(*) begin
    if(when_SramBanks_l75_2) begin
      _zz_sram_2_ports_rsp_valid = 1'b1;
    end else begin
      _zz_sram_2_ports_rsp_valid = 1'b0;
    end
  end

  assign sram_2_ports_rsp_valid = _zz_sram_2_ports_rsp_valid;
  always @(*) begin
    sram_3_ports_rsp_payload_data[63 : 0] = _zz_sram_3_banks_0_bank_port1;
    sram_3_ports_rsp_payload_data[127 : 64] = _zz_sram_3_banks_1_bank_port1;
    sram_3_ports_rsp_payload_data[191 : 128] = _zz_sram_3_banks_2_bank_port1;
    sram_3_ports_rsp_payload_data[255 : 192] = _zz_sram_3_banks_3_bank_port1;
    sram_3_ports_rsp_payload_data[319 : 256] = _zz_sram_3_banks_4_bank_port1;
    sram_3_ports_rsp_payload_data[383 : 320] = _zz_sram_3_banks_5_bank_port1;
    sram_3_ports_rsp_payload_data[447 : 384] = _zz_sram_3_banks_6_bank_port1;
    sram_3_ports_rsp_payload_data[511 : 448] = _zz_sram_3_banks_7_bank_port1;
  end

  assign when_SramBanks_l75_3 = (sram_3_ports_cmd_valid && (sram_3_ports_cmd_payload_wen == 8'h0));
  always @(*) begin
    if(when_SramBanks_l75_3) begin
      _zz_sram_3_ports_rsp_valid = 1'b1;
    end else begin
      _zz_sram_3_ports_rsp_valid = 1'b0;
    end
  end

  assign sram_3_ports_rsp_valid = _zz_sram_3_ports_rsp_valid;

endmodule

module DCache (
  output              stall,
  input               flush,
  input               cpu_cmd_valid,
  output              cpu_cmd_ready,
  input      [63:0]   cpu_cmd_payload_addr,
  input               cpu_cmd_payload_wen,
  input      [63:0]   cpu_cmd_payload_wdata,
  input      [7:0]    cpu_cmd_payload_wstrb,
  input      [2:0]    cpu_cmd_payload_size,
  output              cpu_rsp_valid,
  output     [63:0]   cpu_rsp_payload_data,
  output reg          sram_0_ports_cmd_valid,
  output reg [1:0]    sram_0_ports_cmd_payload_addr,
  output reg [7:0]    sram_0_ports_cmd_payload_wen,
  output reg [511:0]  sram_0_ports_cmd_payload_wdata,
  output reg [63:0]   sram_0_ports_cmd_payload_wstrb,
  input               sram_0_ports_rsp_valid,
  input      [511:0]  sram_0_ports_rsp_payload_data,
  output reg          sram_1_ports_cmd_valid,
  output reg [1:0]    sram_1_ports_cmd_payload_addr,
  output reg [7:0]    sram_1_ports_cmd_payload_wen,
  output reg [511:0]  sram_1_ports_cmd_payload_wdata,
  output reg [63:0]   sram_1_ports_cmd_payload_wstrb,
  input               sram_1_ports_rsp_valid,
  input      [511:0]  sram_1_ports_rsp_payload_data,
  output reg          sram_2_ports_cmd_valid,
  output reg [1:0]    sram_2_ports_cmd_payload_addr,
  output reg [7:0]    sram_2_ports_cmd_payload_wen,
  output reg [511:0]  sram_2_ports_cmd_payload_wdata,
  output reg [63:0]   sram_2_ports_cmd_payload_wstrb,
  input               sram_2_ports_rsp_valid,
  input      [511:0]  sram_2_ports_rsp_payload_data,
  output reg          sram_3_ports_cmd_valid,
  output reg [1:0]    sram_3_ports_cmd_payload_addr,
  output reg [7:0]    sram_3_ports_cmd_payload_wen,
  output reg [511:0]  sram_3_ports_cmd_payload_wdata,
  output reg [63:0]   sram_3_ports_cmd_payload_wstrb,
  input               sram_3_ports_rsp_valid,
  input      [511:0]  sram_3_ports_rsp_payload_data,
  output              next_level_cmd_valid,
  input               next_level_cmd_ready,
  output     [63:0]   next_level_cmd_payload_addr,
  output     [3:0]    next_level_cmd_payload_len,
  output     [2:0]    next_level_cmd_payload_size,
  output              next_level_cmd_payload_wen,
  output     [63:0]   next_level_cmd_payload_wdata,
  output     [7:0]    next_level_cmd_payload_wstrb,
  input               next_level_rsp_valid,
  input      [63:0]   next_level_rsp_payload_data,
  input      [1:0]    next_level_rsp_payload_bresp,
  input               next_level_rsp_payload_rvalid,
  output              cpu_bypass_cmd_valid,
  input               cpu_bypass_cmd_ready,
  output     [63:0]   cpu_bypass_cmd_payload_addr,
  output              cpu_bypass_cmd_payload_wen,
  output     [63:0]   cpu_bypass_cmd_payload_wdata,
  output     [7:0]    cpu_bypass_cmd_payload_wstrb,
  output     [2:0]    cpu_bypass_cmd_payload_size,
  input               cpu_bypass_rsp_valid,
  input      [63:0]   cpu_bypass_rsp_payload_data,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  wire       [63:0]   _zz_bypass_cond_0;
  wire       [31:0]   _zz_bypass_cond_0_1;
  wire       [63:0]   _zz_bypass_cond_0_2;
  wire       [31:0]   _zz_bypass_cond_0_3;
  wire       [63:0]   _zz_bypass_cond_1;
  wire       [31:0]   _zz_bypass_cond_1_1;
  wire       [63:0]   _zz_bypass_cond_1_2;
  wire       [31:0]   _zz_bypass_cond_1_3;
  wire       [63:0]   _zz_bypass_cond_2;
  wire       [31:0]   _zz_bypass_cond_2_1;
  wire       [1:0]    _zz_flush_cnt_valueNext;
  wire       [0:0]    _zz_flush_cnt_valueNext_1;
  wire       [2:0]    _zz_next_level_data_cnt_valueNext;
  wire       [0:0]    _zz_next_level_data_cnt_valueNext_1;
  wire       [6:0]    _zz_next_level_wstrb;
  wire       [7:0]    _zz__zz_cache_hit_gnt_0_3;
  wire       [7:0]    _zz__zz_cache_hit_gnt_0_3_1;
  wire       [3:0]    _zz__zz_cache_hit_gnt_0_3_2;
  wire       [7:0]    _zz__zz_cache_invld_gnt_0_3;
  wire       [7:0]    _zz__zz_cache_invld_gnt_0_3_1;
  wire       [3:0]    _zz__zz_cache_invld_gnt_0_3_2;
  wire       [7:0]    _zz__zz_cache_victim_gnt_0_3;
  wire       [7:0]    _zz__zz_cache_victim_gnt_0_3_1;
  wire       [3:0]    _zz__zz_cache_victim_gnt_0_3_2;
  reg                 _zz__zz_cache_hit_0;
  reg                 _zz__zz_cache_mru_0;
  reg        [55:0]   _zz_cache_tag_0;
  wire       [9:0]    _zz_sram_0_ports_cmd_payload_wdata;
  wire       [9:0]    _zz_sram_0_ports_cmd_payload_wstrb;
  wire       [9:0]    _zz_sram_0_ports_cmd_payload_wstrb_1;
  wire       [3:0]    _zz_sram_0_ports_cmd_payload_wen_1;
  wire       [9:0]    _zz_sram_0_ports_cmd_payload_wdata_1;
  wire       [9:0]    _zz_sram_0_ports_cmd_payload_wstrb_2;
  wire       [9:0]    _zz_sram_0_ports_cmd_payload_wstrb_3;
  reg                 _zz__zz_cache_hit_1;
  reg                 _zz__zz_cache_mru_1;
  reg        [55:0]   _zz_cache_tag_1;
  wire       [9:0]    _zz_sram_1_ports_cmd_payload_wdata;
  wire       [9:0]    _zz_sram_1_ports_cmd_payload_wstrb;
  wire       [9:0]    _zz_sram_1_ports_cmd_payload_wstrb_1;
  wire       [3:0]    _zz_sram_1_ports_cmd_payload_wen_1;
  wire       [9:0]    _zz_sram_1_ports_cmd_payload_wdata_1;
  wire       [9:0]    _zz_sram_1_ports_cmd_payload_wstrb_2;
  wire       [9:0]    _zz_sram_1_ports_cmd_payload_wstrb_3;
  reg                 _zz__zz_cache_hit_2;
  reg                 _zz__zz_cache_mru_2;
  reg        [55:0]   _zz_cache_tag_2;
  wire       [9:0]    _zz_sram_2_ports_cmd_payload_wdata;
  wire       [9:0]    _zz_sram_2_ports_cmd_payload_wstrb;
  wire       [9:0]    _zz_sram_2_ports_cmd_payload_wstrb_1;
  wire       [3:0]    _zz_sram_2_ports_cmd_payload_wen_1;
  wire       [9:0]    _zz_sram_2_ports_cmd_payload_wdata_1;
  wire       [9:0]    _zz_sram_2_ports_cmd_payload_wstrb_2;
  wire       [9:0]    _zz_sram_2_ports_cmd_payload_wstrb_3;
  reg                 _zz__zz_cache_hit_3;
  reg                 _zz__zz_cache_mru_3;
  reg        [55:0]   _zz_cache_tag_3;
  wire       [9:0]    _zz_sram_3_ports_cmd_payload_wdata;
  wire       [9:0]    _zz_sram_3_ports_cmd_payload_wstrb;
  wire       [9:0]    _zz_sram_3_ports_cmd_payload_wstrb_1;
  wire       [3:0]    _zz_sram_3_ports_cmd_payload_wen_1;
  wire       [9:0]    _zz_sram_3_ports_cmd_payload_wdata_1;
  wire       [9:0]    _zz_sram_3_ports_cmd_payload_wstrb_2;
  wire       [9:0]    _zz_sram_3_ports_cmd_payload_wstrb_3;
  reg        [511:0]  _zz__zz_hit_data;
  reg        [63:0]   _zz_hit_data_1;
  reg        [511:0]  _zz__zz_refill_data;
  reg        [63:0]   _zz_refill_data_1;
  reg                 _zz_cpu_rsp_valid;
  reg                 _zz_cpu_rsp_valid_1;
  wire                cpu_stall;
  wire                cpu_bypass_stall;
  reg                 ways_0_metas_0_vld;
  reg        [55:0]   ways_0_metas_0_tag;
  reg                 ways_0_metas_0_mru;
  reg                 ways_0_metas_1_vld;
  reg        [55:0]   ways_0_metas_1_tag;
  reg                 ways_0_metas_1_mru;
  reg                 ways_0_metas_2_vld;
  reg        [55:0]   ways_0_metas_2_tag;
  reg                 ways_0_metas_2_mru;
  reg                 ways_0_metas_3_vld;
  reg        [55:0]   ways_0_metas_3_tag;
  reg                 ways_0_metas_3_mru;
  reg                 ways_1_metas_0_vld;
  reg        [55:0]   ways_1_metas_0_tag;
  reg                 ways_1_metas_0_mru;
  reg                 ways_1_metas_1_vld;
  reg        [55:0]   ways_1_metas_1_tag;
  reg                 ways_1_metas_1_mru;
  reg                 ways_1_metas_2_vld;
  reg        [55:0]   ways_1_metas_2_tag;
  reg                 ways_1_metas_2_mru;
  reg                 ways_1_metas_3_vld;
  reg        [55:0]   ways_1_metas_3_tag;
  reg                 ways_1_metas_3_mru;
  reg                 ways_2_metas_0_vld;
  reg        [55:0]   ways_2_metas_0_tag;
  reg                 ways_2_metas_0_mru;
  reg                 ways_2_metas_1_vld;
  reg        [55:0]   ways_2_metas_1_tag;
  reg                 ways_2_metas_1_mru;
  reg                 ways_2_metas_2_vld;
  reg        [55:0]   ways_2_metas_2_tag;
  reg                 ways_2_metas_2_mru;
  reg                 ways_2_metas_3_vld;
  reg        [55:0]   ways_2_metas_3_tag;
  reg                 ways_2_metas_3_mru;
  reg                 ways_3_metas_0_vld;
  reg        [55:0]   ways_3_metas_0_tag;
  reg                 ways_3_metas_0_mru;
  reg                 ways_3_metas_1_vld;
  reg        [55:0]   ways_3_metas_1_tag;
  reg                 ways_3_metas_1_mru;
  reg                 ways_3_metas_2_vld;
  reg        [55:0]   ways_3_metas_2_tag;
  reg                 ways_3_metas_2_mru;
  reg                 ways_3_metas_3_vld;
  reg        [55:0]   ways_3_metas_3_tag;
  reg                 ways_3_metas_3_mru;
  reg                 cpu_cmd_ready_1;
  wire       [55:0]   cpu_tag;
  wire       [1:0]    cpu_set;
  wire       [1:0]    cpu_bank_addr;
  wire       [2:0]    cpu_bank_index;
  wire                bypass_cond_0;
  wire                bypass_cond_1;
  wire                bypass_cond_2;
  wire                cpu_cmd_fire;
  wire                bypass;
  reg                 bypass_reg;
  reg                 bypass_rsp_valid_d1;
  reg        [63:0]   bypass_rsp_data_d1;
  wire       [55:0]   cache_tag_0;
  wire       [55:0]   cache_tag_1;
  wire       [55:0]   cache_tag_2;
  wire       [55:0]   cache_tag_3;
  wire                cache_hit_0;
  wire                cache_hit_1;
  wire                cache_hit_2;
  wire                cache_hit_3;
  wire                cache_invld_0;
  wire                cache_invld_1;
  wire                cache_invld_2;
  wire                cache_invld_3;
  wire                cache_victim_0;
  wire                cache_victim_1;
  wire                cache_victim_2;
  wire                cache_victim_3;
  wire                cache_mru_0;
  wire                cache_mru_1;
  wire                cache_mru_2;
  wire                cache_mru_3;
  wire                cache_lru_0;
  wire                cache_lru_1;
  wire                cache_lru_2;
  wire                cache_lru_3;
  wire       [1:0]    hit_id;
  wire       [1:0]    evict_id;
  wire       [1:0]    invld_id;
  wire       [1:0]    victim_id;
  wire                mru_full;
  wire                cpu_cmd_fire_1;
  wire                is_hit;
  wire                cpu_cmd_fire_2;
  wire                is_miss;
  wire                is_diff;
  wire                cpu_cmd_fire_3;
  wire                is_write;
  reg                 flush_busy;
  reg                 flush_cnt_willIncrement;
  reg                 flush_cnt_willClear;
  reg        [1:0]    flush_cnt_valueNext;
  reg        [1:0]    flush_cnt_value;
  wire                flush_cnt_willOverflowIfInc;
  wire                flush_cnt_willOverflow;
  wire                flush_done;
  wire                cache_hit_gnt_0;
  wire                cache_hit_gnt_1;
  wire                cache_hit_gnt_2;
  wire                cache_hit_gnt_3;
  wire                cache_victim_gnt_0;
  wire                cache_victim_gnt_1;
  wire                cache_victim_gnt_2;
  wire                cache_victim_gnt_3;
  wire                cache_invld_gnt_0;
  wire                cache_invld_gnt_1;
  wire                cache_invld_gnt_2;
  wire                cache_invld_gnt_3;
  reg        [1:0]    evict_id_miss;
  wire       [511:0]  sram_banks_data_0;
  wire       [511:0]  sram_banks_data_1;
  wire       [511:0]  sram_banks_data_2;
  wire       [511:0]  sram_banks_data_3;
  wire                sram_banks_valid_0;
  wire                sram_banks_valid_1;
  wire                sram_banks_valid_2;
  wire                sram_banks_valid_3;
  reg                 next_level_cmd_valid_1;
  reg                 next_level_data_cnt_willIncrement;
  reg                 next_level_data_cnt_willClear;
  reg        [2:0]    next_level_data_cnt_valueNext;
  reg        [2:0]    next_level_data_cnt_value;
  wire                next_level_data_cnt_willOverflowIfInc;
  wire                next_level_data_cnt_willOverflow;
  wire       [1:0]    next_level_bank_addr;
  wire                next_level_rvalid;
  reg                 next_level_rdone;
  reg                 next_level_wdone;
  wire       [7:0]    next_level_wstrb_tmp;
  wire       [63:0]   next_level_wdata_tmp;
  wire       [7:0]    next_level_wstrb;
  wire       [63:0]   next_level_wdata;
  wire                when_DCache_l145;
  wire                when_DCache_l152;
  wire                when_DCache_l170;
  wire       [3:0]    _zz_cache_hit_gnt_0;
  wire       [3:0]    _zz_cache_hit_gnt_0_1;
  wire       [7:0]    _zz_cache_hit_gnt_0_2;
  wire       [7:0]    _zz_cache_hit_gnt_0_3;
  wire       [3:0]    _zz_cache_hit_gnt_0_4;
  wire       [3:0]    _zz_cache_invld_gnt_0;
  wire       [3:0]    _zz_cache_invld_gnt_0_1;
  wire       [7:0]    _zz_cache_invld_gnt_0_2;
  wire       [7:0]    _zz_cache_invld_gnt_0_3;
  wire       [3:0]    _zz_cache_invld_gnt_0_4;
  wire       [3:0]    _zz_cache_victim_gnt_0;
  wire       [3:0]    _zz_cache_victim_gnt_0_1;
  wire       [7:0]    _zz_cache_victim_gnt_0_2;
  wire       [7:0]    _zz_cache_victim_gnt_0_3;
  wire       [3:0]    _zz_cache_victim_gnt_0_4;
  wire                _zz_hit_id;
  wire                _zz_hit_id_1;
  wire                _zz_invld_id;
  wire                _zz_invld_id_1;
  wire                _zz_victim_id;
  wire                _zz_victim_id_1;
  wire                _zz_cache_hit_0;
  wire                _zz_cache_mru_0;
  wire       [3:0]    _zz_1;
  wire                _zz_2;
  wire                _zz_3;
  wire                _zz_4;
  wire                _zz_5;
  wire                when_DCache_l201;
  reg        [7:0]    _zz_sram_0_ports_cmd_payload_wen;
  wire                when_DCache_l208;
  wire                when_DCache_l215;
  wire       [3:0]    _zz_6;
  wire                _zz_7;
  wire                _zz_8;
  wire                _zz_9;
  wire                _zz_10;
  wire                when_DCache_l237;
  wire                when_DCache_l244;
  wire                when_DCache_l247;
  wire                when_DCache_l252;
  wire                _zz_cache_hit_1;
  wire                _zz_cache_mru_1;
  wire       [3:0]    _zz_11;
  wire                _zz_12;
  wire                _zz_13;
  wire                _zz_14;
  wire                _zz_15;
  wire                when_DCache_l201_1;
  reg        [7:0]    _zz_sram_1_ports_cmd_payload_wen;
  wire                when_DCache_l208_1;
  wire                when_DCache_l215_1;
  wire       [3:0]    _zz_16;
  wire                _zz_17;
  wire                _zz_18;
  wire                _zz_19;
  wire                _zz_20;
  wire                when_DCache_l237_1;
  wire                when_DCache_l244_1;
  wire                when_DCache_l247_1;
  wire                when_DCache_l252_1;
  wire                _zz_cache_hit_2;
  wire                _zz_cache_mru_2;
  wire       [3:0]    _zz_21;
  wire                _zz_22;
  wire                _zz_23;
  wire                _zz_24;
  wire                _zz_25;
  wire                when_DCache_l201_2;
  reg        [7:0]    _zz_sram_2_ports_cmd_payload_wen;
  wire                when_DCache_l208_2;
  wire                when_DCache_l215_2;
  wire       [3:0]    _zz_26;
  wire                _zz_27;
  wire                _zz_28;
  wire                _zz_29;
  wire                _zz_30;
  wire                when_DCache_l237_2;
  wire                when_DCache_l244_2;
  wire                when_DCache_l247_2;
  wire                when_DCache_l252_2;
  wire                _zz_cache_hit_3;
  wire                _zz_cache_mru_3;
  wire       [3:0]    _zz_31;
  wire                _zz_32;
  wire                _zz_33;
  wire                _zz_34;
  wire                _zz_35;
  wire                when_DCache_l201_3;
  reg        [7:0]    _zz_sram_3_ports_cmd_payload_wen;
  wire                when_DCache_l208_3;
  wire                when_DCache_l215_3;
  wire       [3:0]    _zz_36;
  wire                _zz_37;
  wire                _zz_38;
  wire                _zz_39;
  wire                _zz_40;
  wire                when_DCache_l237_3;
  wire                when_DCache_l244_3;
  wire                when_DCache_l247_3;
  wire                when_DCache_l252_3;
  wire                when_DCache_l258;
  wire                when_DCache_l261;
  wire       [511:0]  _zz_hit_data;
  wire       [63:0]   hit_data;
  wire       [511:0]  _zz_refill_data;
  wire       [63:0]   refill_data;
  wire                bypass_stall;
  wire                dcache_stall;
  wire       [63:0]   waddr;
  wire       [63:0]   raddr;
  function [7:0] zz__zz_sram_0_ports_cmd_payload_wen(input dummy);
    begin
      zz__zz_sram_0_ports_cmd_payload_wen = 8'h0;
      zz__zz_sram_0_ports_cmd_payload_wen[0] = 1'b1;
    end
  endfunction
  wire [7:0] _zz_41;
  function [7:0] zz__zz_sram_1_ports_cmd_payload_wen(input dummy);
    begin
      zz__zz_sram_1_ports_cmd_payload_wen = 8'h0;
      zz__zz_sram_1_ports_cmd_payload_wen[0] = 1'b1;
    end
  endfunction
  wire [7:0] _zz_42;
  function [7:0] zz__zz_sram_2_ports_cmd_payload_wen(input dummy);
    begin
      zz__zz_sram_2_ports_cmd_payload_wen = 8'h0;
      zz__zz_sram_2_ports_cmd_payload_wen[0] = 1'b1;
    end
  endfunction
  wire [7:0] _zz_43;
  function [7:0] zz__zz_sram_3_ports_cmd_payload_wen(input dummy);
    begin
      zz__zz_sram_3_ports_cmd_payload_wen = 8'h0;
      zz__zz_sram_3_ports_cmd_payload_wen[0] = 1'b1;
    end
  endfunction
  wire [7:0] _zz_44;

  assign _zz_bypass_cond_0_1 = 32'h10000000;
  assign _zz_bypass_cond_0 = {32'd0, _zz_bypass_cond_0_1};
  assign _zz_bypass_cond_0_3 = 32'h10000fff;
  assign _zz_bypass_cond_0_2 = {32'd0, _zz_bypass_cond_0_3};
  assign _zz_bypass_cond_1_1 = 32'h10001000;
  assign _zz_bypass_cond_1 = {32'd0, _zz_bypass_cond_1_1};
  assign _zz_bypass_cond_1_3 = 32'h10001fff;
  assign _zz_bypass_cond_1_2 = {32'd0, _zz_bypass_cond_1_3};
  assign _zz_bypass_cond_2_1 = 32'h80000000;
  assign _zz_bypass_cond_2 = {32'd0, _zz_bypass_cond_2_1};
  assign _zz_flush_cnt_valueNext_1 = flush_cnt_willIncrement;
  assign _zz_flush_cnt_valueNext = {1'd0, _zz_flush_cnt_valueNext_1};
  assign _zz_next_level_data_cnt_valueNext_1 = next_level_data_cnt_willIncrement;
  assign _zz_next_level_data_cnt_valueNext = {2'd0, _zz_next_level_data_cnt_valueNext_1};
  assign _zz_next_level_wstrb = (7'h0 / 4'b1000);
  assign _zz__zz_cache_hit_gnt_0_3 = (_zz_cache_hit_gnt_0_2 - _zz__zz_cache_hit_gnt_0_3_1);
  assign _zz__zz_cache_hit_gnt_0_3_2 = {_zz_cache_hit_gnt_0[3],{_zz_cache_hit_gnt_0[2],{_zz_cache_hit_gnt_0[1],_zz_cache_hit_gnt_0[0]}}};
  assign _zz__zz_cache_hit_gnt_0_3_1 = {4'd0, _zz__zz_cache_hit_gnt_0_3_2};
  assign _zz__zz_cache_invld_gnt_0_3 = (_zz_cache_invld_gnt_0_2 - _zz__zz_cache_invld_gnt_0_3_1);
  assign _zz__zz_cache_invld_gnt_0_3_2 = {_zz_cache_invld_gnt_0[3],{_zz_cache_invld_gnt_0[2],{_zz_cache_invld_gnt_0[1],_zz_cache_invld_gnt_0[0]}}};
  assign _zz__zz_cache_invld_gnt_0_3_1 = {4'd0, _zz__zz_cache_invld_gnt_0_3_2};
  assign _zz__zz_cache_victim_gnt_0_3 = (_zz_cache_victim_gnt_0_2 - _zz__zz_cache_victim_gnt_0_3_1);
  assign _zz__zz_cache_victim_gnt_0_3_2 = {_zz_cache_victim_gnt_0[3],{_zz_cache_victim_gnt_0[2],{_zz_cache_victim_gnt_0[1],_zz_cache_victim_gnt_0[0]}}};
  assign _zz__zz_cache_victim_gnt_0_3_1 = {4'd0, _zz__zz_cache_victim_gnt_0_3_2};
  assign _zz_sram_0_ports_cmd_payload_wdata = (cpu_bank_index * 7'h40);
  assign _zz_sram_0_ports_cmd_payload_wstrb = (_zz_sram_0_ports_cmd_payload_wstrb_1 / 4'b1000);
  assign _zz_sram_0_ports_cmd_payload_wstrb_1 = (cpu_bank_index * 7'h40);
  assign _zz_sram_0_ports_cmd_payload_wen_1 = (next_level_data_cnt_value * 1'b1);
  assign _zz_sram_0_ports_cmd_payload_wdata_1 = (next_level_data_cnt_value * 7'h40);
  assign _zz_sram_0_ports_cmd_payload_wstrb_2 = (_zz_sram_0_ports_cmd_payload_wstrb_3 / 4'b1000);
  assign _zz_sram_0_ports_cmd_payload_wstrb_3 = (next_level_data_cnt_value * 7'h40);
  assign _zz_sram_1_ports_cmd_payload_wdata = (cpu_bank_index * 7'h40);
  assign _zz_sram_1_ports_cmd_payload_wstrb = (_zz_sram_1_ports_cmd_payload_wstrb_1 / 4'b1000);
  assign _zz_sram_1_ports_cmd_payload_wstrb_1 = (cpu_bank_index * 7'h40);
  assign _zz_sram_1_ports_cmd_payload_wen_1 = (next_level_data_cnt_value * 1'b1);
  assign _zz_sram_1_ports_cmd_payload_wdata_1 = (next_level_data_cnt_value * 7'h40);
  assign _zz_sram_1_ports_cmd_payload_wstrb_2 = (_zz_sram_1_ports_cmd_payload_wstrb_3 / 4'b1000);
  assign _zz_sram_1_ports_cmd_payload_wstrb_3 = (next_level_data_cnt_value * 7'h40);
  assign _zz_sram_2_ports_cmd_payload_wdata = (cpu_bank_index * 7'h40);
  assign _zz_sram_2_ports_cmd_payload_wstrb = (_zz_sram_2_ports_cmd_payload_wstrb_1 / 4'b1000);
  assign _zz_sram_2_ports_cmd_payload_wstrb_1 = (cpu_bank_index * 7'h40);
  assign _zz_sram_2_ports_cmd_payload_wen_1 = (next_level_data_cnt_value * 1'b1);
  assign _zz_sram_2_ports_cmd_payload_wdata_1 = (next_level_data_cnt_value * 7'h40);
  assign _zz_sram_2_ports_cmd_payload_wstrb_2 = (_zz_sram_2_ports_cmd_payload_wstrb_3 / 4'b1000);
  assign _zz_sram_2_ports_cmd_payload_wstrb_3 = (next_level_data_cnt_value * 7'h40);
  assign _zz_sram_3_ports_cmd_payload_wdata = (cpu_bank_index * 7'h40);
  assign _zz_sram_3_ports_cmd_payload_wstrb = (_zz_sram_3_ports_cmd_payload_wstrb_1 / 4'b1000);
  assign _zz_sram_3_ports_cmd_payload_wstrb_1 = (cpu_bank_index * 7'h40);
  assign _zz_sram_3_ports_cmd_payload_wen_1 = (next_level_data_cnt_value * 1'b1);
  assign _zz_sram_3_ports_cmd_payload_wdata_1 = (next_level_data_cnt_value * 7'h40);
  assign _zz_sram_3_ports_cmd_payload_wstrb_2 = (_zz_sram_3_ports_cmd_payload_wstrb_3 / 4'b1000);
  assign _zz_sram_3_ports_cmd_payload_wstrb_3 = (next_level_data_cnt_value * 7'h40);
  always @(*) begin
    case(cpu_set)
      2'b00 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_0_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_0_mru;
        _zz_cache_tag_0 = ways_0_metas_0_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_0_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_0_mru;
        _zz_cache_tag_1 = ways_1_metas_0_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_0_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_0_mru;
        _zz_cache_tag_2 = ways_2_metas_0_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_0_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_0_mru;
        _zz_cache_tag_3 = ways_3_metas_0_tag;
      end
      2'b01 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_1_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_1_mru;
        _zz_cache_tag_0 = ways_0_metas_1_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_1_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_1_mru;
        _zz_cache_tag_1 = ways_1_metas_1_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_1_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_1_mru;
        _zz_cache_tag_2 = ways_2_metas_1_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_1_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_1_mru;
        _zz_cache_tag_3 = ways_3_metas_1_tag;
      end
      2'b10 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_2_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_2_mru;
        _zz_cache_tag_0 = ways_0_metas_2_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_2_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_2_mru;
        _zz_cache_tag_1 = ways_1_metas_2_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_2_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_2_mru;
        _zz_cache_tag_2 = ways_2_metas_2_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_2_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_2_mru;
        _zz_cache_tag_3 = ways_3_metas_2_tag;
      end
      default : begin
        _zz__zz_cache_hit_0 = ways_0_metas_3_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_3_mru;
        _zz_cache_tag_0 = ways_0_metas_3_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_3_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_3_mru;
        _zz_cache_tag_1 = ways_1_metas_3_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_3_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_3_mru;
        _zz_cache_tag_2 = ways_2_metas_3_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_3_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_3_mru;
        _zz_cache_tag_3 = ways_3_metas_3_tag;
      end
    endcase
  end

  always @(*) begin
    case(hit_id)
      2'b00 : begin
        _zz__zz_hit_data = sram_banks_data_0;
        _zz_cpu_rsp_valid = sram_banks_valid_0;
      end
      2'b01 : begin
        _zz__zz_hit_data = sram_banks_data_1;
        _zz_cpu_rsp_valid = sram_banks_valid_1;
      end
      2'b10 : begin
        _zz__zz_hit_data = sram_banks_data_2;
        _zz_cpu_rsp_valid = sram_banks_valid_2;
      end
      default : begin
        _zz__zz_hit_data = sram_banks_data_3;
        _zz_cpu_rsp_valid = sram_banks_valid_3;
      end
    endcase
  end

  always @(*) begin
    case(cpu_bank_index)
      3'b000 : begin
        _zz_hit_data_1 = _zz_hit_data[63 : 0];
        _zz_refill_data_1 = _zz_refill_data[63 : 0];
      end
      3'b001 : begin
        _zz_hit_data_1 = _zz_hit_data[127 : 64];
        _zz_refill_data_1 = _zz_refill_data[127 : 64];
      end
      3'b010 : begin
        _zz_hit_data_1 = _zz_hit_data[191 : 128];
        _zz_refill_data_1 = _zz_refill_data[191 : 128];
      end
      3'b011 : begin
        _zz_hit_data_1 = _zz_hit_data[255 : 192];
        _zz_refill_data_1 = _zz_refill_data[255 : 192];
      end
      3'b100 : begin
        _zz_hit_data_1 = _zz_hit_data[319 : 256];
        _zz_refill_data_1 = _zz_refill_data[319 : 256];
      end
      3'b101 : begin
        _zz_hit_data_1 = _zz_hit_data[383 : 320];
        _zz_refill_data_1 = _zz_refill_data[383 : 320];
      end
      3'b110 : begin
        _zz_hit_data_1 = _zz_hit_data[447 : 384];
        _zz_refill_data_1 = _zz_refill_data[447 : 384];
      end
      default : begin
        _zz_hit_data_1 = _zz_hit_data[511 : 448];
        _zz_refill_data_1 = _zz_refill_data[511 : 448];
      end
    endcase
  end

  always @(*) begin
    case(evict_id_miss)
      2'b00 : begin
        _zz__zz_refill_data = sram_banks_data_0;
        _zz_cpu_rsp_valid_1 = sram_banks_valid_0;
      end
      2'b01 : begin
        _zz__zz_refill_data = sram_banks_data_1;
        _zz_cpu_rsp_valid_1 = sram_banks_valid_1;
      end
      2'b10 : begin
        _zz__zz_refill_data = sram_banks_data_2;
        _zz_cpu_rsp_valid_1 = sram_banks_valid_2;
      end
      default : begin
        _zz__zz_refill_data = sram_banks_data_3;
        _zz_cpu_rsp_valid_1 = sram_banks_valid_3;
      end
    endcase
  end

  assign cpu_tag = cpu_cmd_payload_addr[63 : 8];
  assign cpu_set = cpu_cmd_payload_addr[7 : 6];
  assign cpu_bank_addr = cpu_cmd_payload_addr[7 : 6];
  assign cpu_bank_index = cpu_cmd_payload_addr[5 : 3];
  assign bypass_cond_0 = ((_zz_bypass_cond_0 <= cpu_cmd_payload_addr) && (cpu_cmd_payload_addr <= _zz_bypass_cond_0_2));
  assign bypass_cond_1 = ((_zz_bypass_cond_1 <= cpu_cmd_payload_addr) && (cpu_cmd_payload_addr <= _zz_bypass_cond_1_2));
  assign bypass_cond_2 = (_zz_bypass_cond_2 <= cpu_cmd_payload_addr);
  assign cpu_cmd_fire = (cpu_cmd_valid && cpu_cmd_ready);
  assign bypass = (((bypass_cond_0 || bypass_cond_1) || bypass_cond_2) && cpu_cmd_fire);
  assign cpu_bypass_cmd_valid = bypass;
  assign cpu_bypass_cmd_payload_addr = cpu_cmd_payload_addr;
  assign cpu_bypass_cmd_payload_wen = cpu_cmd_payload_wen;
  assign cpu_bypass_cmd_payload_wdata = cpu_cmd_payload_wdata;
  assign cpu_bypass_cmd_payload_wstrb = cpu_cmd_payload_wstrb;
  assign cpu_bypass_cmd_payload_size = cpu_cmd_payload_size;
  assign mru_full = (&{cache_mru_3,{cache_mru_2,{cache_mru_1,cache_mru_0}}});
  assign cpu_cmd_fire_1 = (cpu_cmd_valid && cpu_cmd_ready);
  assign is_hit = (((|{cache_hit_3,{cache_hit_2,{cache_hit_1,cache_hit_0}}}) && cpu_cmd_fire_1) && (! bypass));
  assign cpu_cmd_fire_2 = (cpu_cmd_valid && cpu_cmd_ready);
  assign is_miss = (((! (|{cache_hit_3,{cache_hit_2,{cache_hit_1,cache_hit_0}}})) && cpu_cmd_fire_2) && (! bypass));
  assign is_diff = (! (|{cache_victim_3,{cache_victim_2,{cache_victim_1,cache_victim_0}}}));
  assign cpu_cmd_fire_3 = (cpu_cmd_valid && cpu_cmd_ready);
  assign is_write = ((cpu_cmd_fire_3 && cpu_cmd_payload_wen) && (! bypass));
  always @(*) begin
    flush_cnt_willIncrement = 1'b0;
    if(!when_DCache_l170) begin
      if(flush_busy) begin
        flush_cnt_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    flush_cnt_willClear = 1'b0;
    if(when_DCache_l170) begin
      flush_cnt_willClear = 1'b1;
    end
  end

  assign flush_cnt_willOverflowIfInc = (flush_cnt_value == 2'b11);
  assign flush_cnt_willOverflow = (flush_cnt_willOverflowIfInc && flush_cnt_willIncrement);
  always @(*) begin
    flush_cnt_valueNext = (flush_cnt_value + _zz_flush_cnt_valueNext);
    if(flush_cnt_willClear) begin
      flush_cnt_valueNext = 2'b00;
    end
  end

  assign flush_done = (flush_busy && (flush_cnt_value == 2'b11));
  always @(*) begin
    next_level_data_cnt_willIncrement = 1'b0;
    if(!when_DCache_l152) begin
      if(!next_level_rdone) begin
        if(next_level_rvalid) begin
          next_level_data_cnt_willIncrement = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    next_level_data_cnt_willClear = 1'b0;
    if(when_DCache_l152) begin
      next_level_data_cnt_willClear = 1'b1;
    end else begin
      if(next_level_rdone) begin
        next_level_data_cnt_willClear = 1'b1;
      end
    end
  end

  assign next_level_data_cnt_willOverflowIfInc = (next_level_data_cnt_value == 3'b111);
  assign next_level_data_cnt_willOverflow = (next_level_data_cnt_willOverflowIfInc && next_level_data_cnt_willIncrement);
  always @(*) begin
    next_level_data_cnt_valueNext = (next_level_data_cnt_value + _zz_next_level_data_cnt_valueNext);
    if(next_level_data_cnt_willClear) begin
      next_level_data_cnt_valueNext = 3'b000;
    end
  end

  assign next_level_bank_addr = cpu_cmd_payload_addr[7 : 6];
  assign next_level_rvalid = (next_level_rsp_valid && next_level_rsp_payload_rvalid);
  assign next_level_wstrb_tmp = cpu_cmd_payload_wstrb;
  assign next_level_wdata_tmp = cpu_cmd_payload_wdata;
  assign next_level_wstrb = (next_level_wstrb_tmp <<< _zz_next_level_wstrb);
  assign next_level_wdata = (next_level_wdata_tmp <<< 7'h0);
  assign when_DCache_l145 = (is_miss || is_write);
  assign when_DCache_l152 = (is_miss && (! is_write));
  assign when_DCache_l170 = (flush_busy && (flush_cnt_value == 2'b11));
  assign _zz_cache_hit_gnt_0 = 4'b0001;
  assign _zz_cache_hit_gnt_0_1 = {cache_hit_3,{cache_hit_2,{cache_hit_1,cache_hit_0}}};
  assign _zz_cache_hit_gnt_0_2 = {_zz_cache_hit_gnt_0_1,_zz_cache_hit_gnt_0_1};
  assign _zz_cache_hit_gnt_0_3 = (_zz_cache_hit_gnt_0_2 & (~ _zz__zz_cache_hit_gnt_0_3));
  assign _zz_cache_hit_gnt_0_4 = (_zz_cache_hit_gnt_0_3[7 : 4] | _zz_cache_hit_gnt_0_3[3 : 0]);
  assign cache_hit_gnt_0 = _zz_cache_hit_gnt_0_4[0];
  assign cache_hit_gnt_1 = _zz_cache_hit_gnt_0_4[1];
  assign cache_hit_gnt_2 = _zz_cache_hit_gnt_0_4[2];
  assign cache_hit_gnt_3 = _zz_cache_hit_gnt_0_4[3];
  assign _zz_cache_invld_gnt_0 = 4'b0001;
  assign _zz_cache_invld_gnt_0_1 = {cache_invld_3,{cache_invld_2,{cache_invld_1,cache_invld_0}}};
  assign _zz_cache_invld_gnt_0_2 = {_zz_cache_invld_gnt_0_1,_zz_cache_invld_gnt_0_1};
  assign _zz_cache_invld_gnt_0_3 = (_zz_cache_invld_gnt_0_2 & (~ _zz__zz_cache_invld_gnt_0_3));
  assign _zz_cache_invld_gnt_0_4 = (_zz_cache_invld_gnt_0_3[7 : 4] | _zz_cache_invld_gnt_0_3[3 : 0]);
  assign cache_invld_gnt_0 = _zz_cache_invld_gnt_0_4[0];
  assign cache_invld_gnt_1 = _zz_cache_invld_gnt_0_4[1];
  assign cache_invld_gnt_2 = _zz_cache_invld_gnt_0_4[2];
  assign cache_invld_gnt_3 = _zz_cache_invld_gnt_0_4[3];
  assign _zz_cache_victim_gnt_0 = 4'b0001;
  assign _zz_cache_victim_gnt_0_1 = {cache_victim_3,{cache_victim_2,{cache_victim_1,cache_victim_0}}};
  assign _zz_cache_victim_gnt_0_2 = {_zz_cache_victim_gnt_0_1,_zz_cache_victim_gnt_0_1};
  assign _zz_cache_victim_gnt_0_3 = (_zz_cache_victim_gnt_0_2 & (~ _zz__zz_cache_victim_gnt_0_3));
  assign _zz_cache_victim_gnt_0_4 = (_zz_cache_victim_gnt_0_3[7 : 4] | _zz_cache_victim_gnt_0_3[3 : 0]);
  assign cache_victim_gnt_0 = _zz_cache_victim_gnt_0_4[0];
  assign cache_victim_gnt_1 = _zz_cache_victim_gnt_0_4[1];
  assign cache_victim_gnt_2 = _zz_cache_victim_gnt_0_4[2];
  assign cache_victim_gnt_3 = _zz_cache_victim_gnt_0_4[3];
  assign _zz_hit_id = (cache_hit_gnt_1 || cache_hit_gnt_3);
  assign _zz_hit_id_1 = (cache_hit_gnt_2 || cache_hit_gnt_3);
  assign hit_id = {_zz_hit_id_1,_zz_hit_id};
  assign _zz_invld_id = (cache_invld_gnt_1 || cache_invld_gnt_3);
  assign _zz_invld_id_1 = (cache_invld_gnt_2 || cache_invld_gnt_3);
  assign invld_id = {_zz_invld_id_1,_zz_invld_id};
  assign _zz_victim_id = (cache_victim_gnt_1 || cache_victim_gnt_3);
  assign _zz_victim_id_1 = (cache_victim_gnt_2 || cache_victim_gnt_3);
  assign victim_id = {_zz_victim_id_1,_zz_victim_id};
  assign evict_id = (is_diff ? invld_id : victim_id);
  assign _zz_cache_hit_0 = _zz__zz_cache_hit_0;
  assign _zz_cache_mru_0 = _zz__zz_cache_mru_0;
  assign _zz_1 = ({3'd0,1'b1} <<< cpu_set);
  assign _zz_2 = _zz_1[0];
  assign _zz_3 = _zz_1[1];
  assign _zz_4 = _zz_1[2];
  assign _zz_5 = _zz_1[3];
  assign cache_tag_0 = _zz_cache_tag_0;
  assign cache_hit_0 = ((cache_tag_0 == cpu_tag) && _zz_cache_hit_0);
  assign cache_mru_0 = _zz_cache_mru_0;
  assign cache_invld_0 = (! _zz_cache_hit_0);
  assign cache_lru_0 = (! _zz_cache_mru_0);
  assign cache_victim_0 = (cache_invld_0 && cache_lru_0);
  assign sram_banks_data_0 = sram_0_ports_rsp_payload_data;
  assign sram_banks_valid_0 = sram_0_ports_rsp_valid;
  assign when_DCache_l201 = (is_hit && (2'b00 == hit_id));
  always @(*) begin
    if(when_DCache_l201) begin
      sram_0_ports_cmd_payload_addr = cpu_bank_addr;
    end else begin
      if(when_DCache_l208) begin
        sram_0_ports_cmd_payload_addr = cpu_bank_addr;
      end else begin
        if(when_DCache_l215) begin
          sram_0_ports_cmd_payload_addr = next_level_bank_addr;
        end else begin
          sram_0_ports_cmd_payload_addr = 2'b00;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l201) begin
      sram_0_ports_cmd_valid = 1'b1;
    end else begin
      if(when_DCache_l208) begin
        sram_0_ports_cmd_valid = 1'b1;
      end else begin
        if(when_DCache_l215) begin
          sram_0_ports_cmd_valid = 1'b1;
        end else begin
          sram_0_ports_cmd_valid = 1'b0;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l201) begin
      sram_0_ports_cmd_payload_wen = ({7'h0,cpu_cmd_payload_wen} <<< cpu_bank_index);
    end else begin
      if(when_DCache_l208) begin
        sram_0_ports_cmd_payload_wen = 8'h0;
      end else begin
        if(when_DCache_l215) begin
          sram_0_ports_cmd_payload_wen = (_zz_sram_0_ports_cmd_payload_wen <<< _zz_sram_0_ports_cmd_payload_wen_1);
        end else begin
          sram_0_ports_cmd_payload_wen = 8'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l201) begin
      sram_0_ports_cmd_payload_wdata = ({448'h0,cpu_cmd_payload_wdata} <<< _zz_sram_0_ports_cmd_payload_wdata);
    end else begin
      if(when_DCache_l208) begin
        sram_0_ports_cmd_payload_wdata = 512'h0;
      end else begin
        if(when_DCache_l215) begin
          sram_0_ports_cmd_payload_wdata = ({448'h0,next_level_rsp_payload_data} <<< _zz_sram_0_ports_cmd_payload_wdata_1);
        end else begin
          sram_0_ports_cmd_payload_wdata = 512'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l201) begin
      sram_0_ports_cmd_payload_wstrb = ({56'h0,cpu_cmd_payload_wstrb} <<< _zz_sram_0_ports_cmd_payload_wstrb);
    end else begin
      if(when_DCache_l208) begin
        sram_0_ports_cmd_payload_wstrb = 64'h0;
      end else begin
        if(when_DCache_l215) begin
          sram_0_ports_cmd_payload_wstrb = ({56'h0,8'hff} <<< _zz_sram_0_ports_cmd_payload_wstrb_2);
        end else begin
          sram_0_ports_cmd_payload_wstrb = 64'h0;
        end
      end
    end
  end

  assign _zz_41 = zz__zz_sram_0_ports_cmd_payload_wen(1'b0);
  always @(*) _zz_sram_0_ports_cmd_payload_wen = _zz_41;
  assign when_DCache_l208 = ((next_level_rdone && (! is_write)) && (2'b00 == evict_id_miss));
  assign when_DCache_l215 = (next_level_rvalid && (2'b00 == evict_id_miss));
  assign _zz_6 = ({3'd0,1'b1} <<< flush_cnt_value);
  assign _zz_7 = _zz_6[0];
  assign _zz_8 = _zz_6[1];
  assign _zz_9 = _zz_6[2];
  assign _zz_10 = _zz_6[3];
  assign when_DCache_l237 = (is_hit && mru_full);
  assign when_DCache_l244 = (is_hit && cache_hit_0);
  assign when_DCache_l247 = (next_level_rdone && (2'b00 == evict_id_miss));
  assign when_DCache_l252 = (next_level_rdone && (2'b00 == evict_id_miss));
  assign _zz_cache_hit_1 = _zz__zz_cache_hit_1;
  assign _zz_cache_mru_1 = _zz__zz_cache_mru_1;
  assign _zz_11 = ({3'd0,1'b1} <<< cpu_set);
  assign _zz_12 = _zz_11[0];
  assign _zz_13 = _zz_11[1];
  assign _zz_14 = _zz_11[2];
  assign _zz_15 = _zz_11[3];
  assign cache_tag_1 = _zz_cache_tag_1;
  assign cache_hit_1 = ((cache_tag_1 == cpu_tag) && _zz_cache_hit_1);
  assign cache_mru_1 = _zz_cache_mru_1;
  assign cache_invld_1 = (! _zz_cache_hit_1);
  assign cache_lru_1 = (! _zz_cache_mru_1);
  assign cache_victim_1 = (cache_invld_1 && cache_lru_1);
  assign sram_banks_data_1 = sram_1_ports_rsp_payload_data;
  assign sram_banks_valid_1 = sram_1_ports_rsp_valid;
  assign when_DCache_l201_1 = (is_hit && (2'b01 == hit_id));
  always @(*) begin
    if(when_DCache_l201_1) begin
      sram_1_ports_cmd_payload_addr = cpu_bank_addr;
    end else begin
      if(when_DCache_l208_1) begin
        sram_1_ports_cmd_payload_addr = cpu_bank_addr;
      end else begin
        if(when_DCache_l215_1) begin
          sram_1_ports_cmd_payload_addr = next_level_bank_addr;
        end else begin
          sram_1_ports_cmd_payload_addr = 2'b00;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l201_1) begin
      sram_1_ports_cmd_valid = 1'b1;
    end else begin
      if(when_DCache_l208_1) begin
        sram_1_ports_cmd_valid = 1'b1;
      end else begin
        if(when_DCache_l215_1) begin
          sram_1_ports_cmd_valid = 1'b1;
        end else begin
          sram_1_ports_cmd_valid = 1'b0;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l201_1) begin
      sram_1_ports_cmd_payload_wen = ({7'h0,cpu_cmd_payload_wen} <<< cpu_bank_index);
    end else begin
      if(when_DCache_l208_1) begin
        sram_1_ports_cmd_payload_wen = 8'h0;
      end else begin
        if(when_DCache_l215_1) begin
          sram_1_ports_cmd_payload_wen = (_zz_sram_1_ports_cmd_payload_wen <<< _zz_sram_1_ports_cmd_payload_wen_1);
        end else begin
          sram_1_ports_cmd_payload_wen = 8'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l201_1) begin
      sram_1_ports_cmd_payload_wdata = ({448'h0,cpu_cmd_payload_wdata} <<< _zz_sram_1_ports_cmd_payload_wdata);
    end else begin
      if(when_DCache_l208_1) begin
        sram_1_ports_cmd_payload_wdata = 512'h0;
      end else begin
        if(when_DCache_l215_1) begin
          sram_1_ports_cmd_payload_wdata = ({448'h0,next_level_rsp_payload_data} <<< _zz_sram_1_ports_cmd_payload_wdata_1);
        end else begin
          sram_1_ports_cmd_payload_wdata = 512'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l201_1) begin
      sram_1_ports_cmd_payload_wstrb = ({56'h0,cpu_cmd_payload_wstrb} <<< _zz_sram_1_ports_cmd_payload_wstrb);
    end else begin
      if(when_DCache_l208_1) begin
        sram_1_ports_cmd_payload_wstrb = 64'h0;
      end else begin
        if(when_DCache_l215_1) begin
          sram_1_ports_cmd_payload_wstrb = ({56'h0,8'hff} <<< _zz_sram_1_ports_cmd_payload_wstrb_2);
        end else begin
          sram_1_ports_cmd_payload_wstrb = 64'h0;
        end
      end
    end
  end

  assign _zz_42 = zz__zz_sram_1_ports_cmd_payload_wen(1'b0);
  always @(*) _zz_sram_1_ports_cmd_payload_wen = _zz_42;
  assign when_DCache_l208_1 = ((next_level_rdone && (! is_write)) && (2'b01 == evict_id_miss));
  assign when_DCache_l215_1 = (next_level_rvalid && (2'b01 == evict_id_miss));
  assign _zz_16 = ({3'd0,1'b1} <<< flush_cnt_value);
  assign _zz_17 = _zz_16[0];
  assign _zz_18 = _zz_16[1];
  assign _zz_19 = _zz_16[2];
  assign _zz_20 = _zz_16[3];
  assign when_DCache_l237_1 = (is_hit && mru_full);
  assign when_DCache_l244_1 = (is_hit && cache_hit_1);
  assign when_DCache_l247_1 = (next_level_rdone && (2'b01 == evict_id_miss));
  assign when_DCache_l252_1 = (next_level_rdone && (2'b01 == evict_id_miss));
  assign _zz_cache_hit_2 = _zz__zz_cache_hit_2;
  assign _zz_cache_mru_2 = _zz__zz_cache_mru_2;
  assign _zz_21 = ({3'd0,1'b1} <<< cpu_set);
  assign _zz_22 = _zz_21[0];
  assign _zz_23 = _zz_21[1];
  assign _zz_24 = _zz_21[2];
  assign _zz_25 = _zz_21[3];
  assign cache_tag_2 = _zz_cache_tag_2;
  assign cache_hit_2 = ((cache_tag_2 == cpu_tag) && _zz_cache_hit_2);
  assign cache_mru_2 = _zz_cache_mru_2;
  assign cache_invld_2 = (! _zz_cache_hit_2);
  assign cache_lru_2 = (! _zz_cache_mru_2);
  assign cache_victim_2 = (cache_invld_2 && cache_lru_2);
  assign sram_banks_data_2 = sram_2_ports_rsp_payload_data;
  assign sram_banks_valid_2 = sram_2_ports_rsp_valid;
  assign when_DCache_l201_2 = (is_hit && (2'b10 == hit_id));
  always @(*) begin
    if(when_DCache_l201_2) begin
      sram_2_ports_cmd_payload_addr = cpu_bank_addr;
    end else begin
      if(when_DCache_l208_2) begin
        sram_2_ports_cmd_payload_addr = cpu_bank_addr;
      end else begin
        if(when_DCache_l215_2) begin
          sram_2_ports_cmd_payload_addr = next_level_bank_addr;
        end else begin
          sram_2_ports_cmd_payload_addr = 2'b00;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l201_2) begin
      sram_2_ports_cmd_valid = 1'b1;
    end else begin
      if(when_DCache_l208_2) begin
        sram_2_ports_cmd_valid = 1'b1;
      end else begin
        if(when_DCache_l215_2) begin
          sram_2_ports_cmd_valid = 1'b1;
        end else begin
          sram_2_ports_cmd_valid = 1'b0;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l201_2) begin
      sram_2_ports_cmd_payload_wen = ({7'h0,cpu_cmd_payload_wen} <<< cpu_bank_index);
    end else begin
      if(when_DCache_l208_2) begin
        sram_2_ports_cmd_payload_wen = 8'h0;
      end else begin
        if(when_DCache_l215_2) begin
          sram_2_ports_cmd_payload_wen = (_zz_sram_2_ports_cmd_payload_wen <<< _zz_sram_2_ports_cmd_payload_wen_1);
        end else begin
          sram_2_ports_cmd_payload_wen = 8'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l201_2) begin
      sram_2_ports_cmd_payload_wdata = ({448'h0,cpu_cmd_payload_wdata} <<< _zz_sram_2_ports_cmd_payload_wdata);
    end else begin
      if(when_DCache_l208_2) begin
        sram_2_ports_cmd_payload_wdata = 512'h0;
      end else begin
        if(when_DCache_l215_2) begin
          sram_2_ports_cmd_payload_wdata = ({448'h0,next_level_rsp_payload_data} <<< _zz_sram_2_ports_cmd_payload_wdata_1);
        end else begin
          sram_2_ports_cmd_payload_wdata = 512'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l201_2) begin
      sram_2_ports_cmd_payload_wstrb = ({56'h0,cpu_cmd_payload_wstrb} <<< _zz_sram_2_ports_cmd_payload_wstrb);
    end else begin
      if(when_DCache_l208_2) begin
        sram_2_ports_cmd_payload_wstrb = 64'h0;
      end else begin
        if(when_DCache_l215_2) begin
          sram_2_ports_cmd_payload_wstrb = ({56'h0,8'hff} <<< _zz_sram_2_ports_cmd_payload_wstrb_2);
        end else begin
          sram_2_ports_cmd_payload_wstrb = 64'h0;
        end
      end
    end
  end

  assign _zz_43 = zz__zz_sram_2_ports_cmd_payload_wen(1'b0);
  always @(*) _zz_sram_2_ports_cmd_payload_wen = _zz_43;
  assign when_DCache_l208_2 = ((next_level_rdone && (! is_write)) && (2'b10 == evict_id_miss));
  assign when_DCache_l215_2 = (next_level_rvalid && (2'b10 == evict_id_miss));
  assign _zz_26 = ({3'd0,1'b1} <<< flush_cnt_value);
  assign _zz_27 = _zz_26[0];
  assign _zz_28 = _zz_26[1];
  assign _zz_29 = _zz_26[2];
  assign _zz_30 = _zz_26[3];
  assign when_DCache_l237_2 = (is_hit && mru_full);
  assign when_DCache_l244_2 = (is_hit && cache_hit_2);
  assign when_DCache_l247_2 = (next_level_rdone && (2'b10 == evict_id_miss));
  assign when_DCache_l252_2 = (next_level_rdone && (2'b10 == evict_id_miss));
  assign _zz_cache_hit_3 = _zz__zz_cache_hit_3;
  assign _zz_cache_mru_3 = _zz__zz_cache_mru_3;
  assign _zz_31 = ({3'd0,1'b1} <<< cpu_set);
  assign _zz_32 = _zz_31[0];
  assign _zz_33 = _zz_31[1];
  assign _zz_34 = _zz_31[2];
  assign _zz_35 = _zz_31[3];
  assign cache_tag_3 = _zz_cache_tag_3;
  assign cache_hit_3 = ((cache_tag_3 == cpu_tag) && _zz_cache_hit_3);
  assign cache_mru_3 = _zz_cache_mru_3;
  assign cache_invld_3 = (! _zz_cache_hit_3);
  assign cache_lru_3 = (! _zz_cache_mru_3);
  assign cache_victim_3 = (cache_invld_3 && cache_lru_3);
  assign sram_banks_data_3 = sram_3_ports_rsp_payload_data;
  assign sram_banks_valid_3 = sram_3_ports_rsp_valid;
  assign when_DCache_l201_3 = (is_hit && (2'b11 == hit_id));
  always @(*) begin
    if(when_DCache_l201_3) begin
      sram_3_ports_cmd_payload_addr = cpu_bank_addr;
    end else begin
      if(when_DCache_l208_3) begin
        sram_3_ports_cmd_payload_addr = cpu_bank_addr;
      end else begin
        if(when_DCache_l215_3) begin
          sram_3_ports_cmd_payload_addr = next_level_bank_addr;
        end else begin
          sram_3_ports_cmd_payload_addr = 2'b00;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l201_3) begin
      sram_3_ports_cmd_valid = 1'b1;
    end else begin
      if(when_DCache_l208_3) begin
        sram_3_ports_cmd_valid = 1'b1;
      end else begin
        if(when_DCache_l215_3) begin
          sram_3_ports_cmd_valid = 1'b1;
        end else begin
          sram_3_ports_cmd_valid = 1'b0;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l201_3) begin
      sram_3_ports_cmd_payload_wen = ({7'h0,cpu_cmd_payload_wen} <<< cpu_bank_index);
    end else begin
      if(when_DCache_l208_3) begin
        sram_3_ports_cmd_payload_wen = 8'h0;
      end else begin
        if(when_DCache_l215_3) begin
          sram_3_ports_cmd_payload_wen = (_zz_sram_3_ports_cmd_payload_wen <<< _zz_sram_3_ports_cmd_payload_wen_1);
        end else begin
          sram_3_ports_cmd_payload_wen = 8'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l201_3) begin
      sram_3_ports_cmd_payload_wdata = ({448'h0,cpu_cmd_payload_wdata} <<< _zz_sram_3_ports_cmd_payload_wdata);
    end else begin
      if(when_DCache_l208_3) begin
        sram_3_ports_cmd_payload_wdata = 512'h0;
      end else begin
        if(when_DCache_l215_3) begin
          sram_3_ports_cmd_payload_wdata = ({448'h0,next_level_rsp_payload_data} <<< _zz_sram_3_ports_cmd_payload_wdata_1);
        end else begin
          sram_3_ports_cmd_payload_wdata = 512'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l201_3) begin
      sram_3_ports_cmd_payload_wstrb = ({56'h0,cpu_cmd_payload_wstrb} <<< _zz_sram_3_ports_cmd_payload_wstrb);
    end else begin
      if(when_DCache_l208_3) begin
        sram_3_ports_cmd_payload_wstrb = 64'h0;
      end else begin
        if(when_DCache_l215_3) begin
          sram_3_ports_cmd_payload_wstrb = ({56'h0,8'hff} <<< _zz_sram_3_ports_cmd_payload_wstrb_2);
        end else begin
          sram_3_ports_cmd_payload_wstrb = 64'h0;
        end
      end
    end
  end

  assign _zz_44 = zz__zz_sram_3_ports_cmd_payload_wen(1'b0);
  always @(*) _zz_sram_3_ports_cmd_payload_wen = _zz_44;
  assign when_DCache_l208_3 = ((next_level_rdone && (! is_write)) && (2'b11 == evict_id_miss));
  assign when_DCache_l215_3 = (next_level_rvalid && (2'b11 == evict_id_miss));
  assign _zz_36 = ({3'd0,1'b1} <<< flush_cnt_value);
  assign _zz_37 = _zz_36[0];
  assign _zz_38 = _zz_36[1];
  assign _zz_39 = _zz_36[2];
  assign _zz_40 = _zz_36[3];
  assign when_DCache_l237_3 = (is_hit && mru_full);
  assign when_DCache_l244_3 = (is_hit && cache_hit_3);
  assign when_DCache_l247_3 = (next_level_rdone && (2'b11 == evict_id_miss));
  assign when_DCache_l252_3 = (next_level_rdone && (2'b11 == evict_id_miss));
  assign when_DCache_l258 = (((flush || is_miss) || is_write) || bypass);
  assign when_DCache_l261 = (((flush_done || next_level_rdone) || next_level_wdone) || bypass_rsp_valid_d1);
  assign _zz_hit_data = _zz__zz_hit_data;
  assign hit_data = _zz_hit_data_1;
  assign _zz_refill_data = _zz__zz_refill_data;
  assign refill_data = _zz_refill_data_1;
  assign cpu_rsp_payload_data = (bypass_reg ? bypass_rsp_data_d1 : (is_hit ? hit_data : refill_data));
  assign cpu_rsp_valid = (bypass_reg ? bypass_rsp_valid_d1 : (is_hit ? _zz_cpu_rsp_valid : _zz_cpu_rsp_valid_1));
  assign cpu_cmd_ready = cpu_cmd_ready_1;
  assign bypass_stall = (((! cpu_cmd_ready) && (! bypass_rsp_valid_d1)) || bypass);
  assign dcache_stall = (((is_miss || is_write) || bypass_stall) && (! next_level_wdone));
  assign stall = dcache_stall;
  assign waddr = {cpu_cmd_payload_addr[63 : 3],3'b000};
  assign raddr = {cpu_cmd_payload_addr[63 : 6],6'h0};
  assign next_level_cmd_payload_addr = (cpu_cmd_payload_wen ? waddr : raddr);
  assign next_level_cmd_payload_len = (cpu_cmd_payload_wen ? 4'b0000 : 4'b0111);
  assign next_level_cmd_payload_size = 3'b011;
  assign next_level_cmd_payload_wen = cpu_cmd_payload_wen;
  assign next_level_cmd_payload_wdata = next_level_wdata;
  assign next_level_cmd_payload_wstrb = next_level_wstrb;
  assign next_level_cmd_valid = next_level_cmd_valid_1;
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      ways_0_metas_0_vld <= 1'b0;
      ways_0_metas_0_tag <= 56'h0;
      ways_0_metas_0_mru <= 1'b0;
      ways_0_metas_1_vld <= 1'b0;
      ways_0_metas_1_tag <= 56'h0;
      ways_0_metas_1_mru <= 1'b0;
      ways_0_metas_2_vld <= 1'b0;
      ways_0_metas_2_tag <= 56'h0;
      ways_0_metas_2_mru <= 1'b0;
      ways_0_metas_3_vld <= 1'b0;
      ways_0_metas_3_tag <= 56'h0;
      ways_0_metas_3_mru <= 1'b0;
      ways_1_metas_0_vld <= 1'b0;
      ways_1_metas_0_tag <= 56'h0;
      ways_1_metas_0_mru <= 1'b0;
      ways_1_metas_1_vld <= 1'b0;
      ways_1_metas_1_tag <= 56'h0;
      ways_1_metas_1_mru <= 1'b0;
      ways_1_metas_2_vld <= 1'b0;
      ways_1_metas_2_tag <= 56'h0;
      ways_1_metas_2_mru <= 1'b0;
      ways_1_metas_3_vld <= 1'b0;
      ways_1_metas_3_tag <= 56'h0;
      ways_1_metas_3_mru <= 1'b0;
      ways_2_metas_0_vld <= 1'b0;
      ways_2_metas_0_tag <= 56'h0;
      ways_2_metas_0_mru <= 1'b0;
      ways_2_metas_1_vld <= 1'b0;
      ways_2_metas_1_tag <= 56'h0;
      ways_2_metas_1_mru <= 1'b0;
      ways_2_metas_2_vld <= 1'b0;
      ways_2_metas_2_tag <= 56'h0;
      ways_2_metas_2_mru <= 1'b0;
      ways_2_metas_3_vld <= 1'b0;
      ways_2_metas_3_tag <= 56'h0;
      ways_2_metas_3_mru <= 1'b0;
      ways_3_metas_0_vld <= 1'b0;
      ways_3_metas_0_tag <= 56'h0;
      ways_3_metas_0_mru <= 1'b0;
      ways_3_metas_1_vld <= 1'b0;
      ways_3_metas_1_tag <= 56'h0;
      ways_3_metas_1_mru <= 1'b0;
      ways_3_metas_2_vld <= 1'b0;
      ways_3_metas_2_tag <= 56'h0;
      ways_3_metas_2_mru <= 1'b0;
      ways_3_metas_3_vld <= 1'b0;
      ways_3_metas_3_tag <= 56'h0;
      ways_3_metas_3_mru <= 1'b0;
      cpu_cmd_ready_1 <= 1'b1;
      bypass_reg <= 1'b0;
      flush_busy <= 1'b0;
      flush_cnt_value <= 2'b00;
      next_level_cmd_valid_1 <= 1'b0;
      next_level_data_cnt_value <= 3'b000;
    end else begin
      if(bypass) begin
        bypass_reg <= 1'b1;
      end else begin
        if(bypass_rsp_valid_d1) begin
          bypass_reg <= 1'b0;
        end
      end
      flush_cnt_value <= flush_cnt_valueNext;
      next_level_data_cnt_value <= next_level_data_cnt_valueNext;
      if(when_DCache_l145) begin
        next_level_cmd_valid_1 <= 1'b1;
      end else begin
        next_level_cmd_valid_1 <= 1'b0;
      end
      if(flush) begin
        flush_busy <= 1'b1;
      end else begin
        if(flush_done) begin
          flush_busy <= 1'b0;
        end
      end
      if(flush_busy) begin
        if(_zz_7) begin
          ways_0_metas_0_mru <= 1'b0;
        end
        if(_zz_8) begin
          ways_0_metas_1_mru <= 1'b0;
        end
        if(_zz_9) begin
          ways_0_metas_2_mru <= 1'b0;
        end
        if(_zz_10) begin
          ways_0_metas_3_mru <= 1'b0;
        end
        if(_zz_7) begin
          ways_0_metas_0_vld <= 1'b0;
        end
        if(_zz_8) begin
          ways_0_metas_1_vld <= 1'b0;
        end
        if(_zz_9) begin
          ways_0_metas_2_vld <= 1'b0;
        end
        if(_zz_10) begin
          ways_0_metas_3_vld <= 1'b0;
        end
      end else begin
        if(when_DCache_l237) begin
          if(cache_hit_0) begin
            if(_zz_2) begin
              ways_0_metas_0_mru <= 1'b1;
            end
            if(_zz_3) begin
              ways_0_metas_1_mru <= 1'b1;
            end
            if(_zz_4) begin
              ways_0_metas_2_mru <= 1'b1;
            end
            if(_zz_5) begin
              ways_0_metas_3_mru <= 1'b1;
            end
          end else begin
            if(_zz_2) begin
              ways_0_metas_0_mru <= 1'b0;
            end
            if(_zz_3) begin
              ways_0_metas_1_mru <= 1'b0;
            end
            if(_zz_4) begin
              ways_0_metas_2_mru <= 1'b0;
            end
            if(_zz_5) begin
              ways_0_metas_3_mru <= 1'b0;
            end
          end
        end else begin
          if(when_DCache_l244) begin
            if(_zz_2) begin
              ways_0_metas_0_mru <= 1'b1;
            end
            if(_zz_3) begin
              ways_0_metas_1_mru <= 1'b1;
            end
            if(_zz_4) begin
              ways_0_metas_2_mru <= 1'b1;
            end
            if(_zz_5) begin
              ways_0_metas_3_mru <= 1'b1;
            end
          end else begin
            if(when_DCache_l247) begin
              if(_zz_2) begin
                ways_0_metas_0_vld <= 1'b1;
              end
              if(_zz_3) begin
                ways_0_metas_1_vld <= 1'b1;
              end
              if(_zz_4) begin
                ways_0_metas_2_vld <= 1'b1;
              end
              if(_zz_5) begin
                ways_0_metas_3_vld <= 1'b1;
              end
            end
          end
        end
      end
      if(when_DCache_l252) begin
        if(_zz_2) begin
          ways_0_metas_0_tag <= cpu_tag;
        end
        if(_zz_3) begin
          ways_0_metas_1_tag <= cpu_tag;
        end
        if(_zz_4) begin
          ways_0_metas_2_tag <= cpu_tag;
        end
        if(_zz_5) begin
          ways_0_metas_3_tag <= cpu_tag;
        end
      end
      if(flush_busy) begin
        if(_zz_17) begin
          ways_1_metas_0_mru <= 1'b0;
        end
        if(_zz_18) begin
          ways_1_metas_1_mru <= 1'b0;
        end
        if(_zz_19) begin
          ways_1_metas_2_mru <= 1'b0;
        end
        if(_zz_20) begin
          ways_1_metas_3_mru <= 1'b0;
        end
        if(_zz_17) begin
          ways_1_metas_0_vld <= 1'b0;
        end
        if(_zz_18) begin
          ways_1_metas_1_vld <= 1'b0;
        end
        if(_zz_19) begin
          ways_1_metas_2_vld <= 1'b0;
        end
        if(_zz_20) begin
          ways_1_metas_3_vld <= 1'b0;
        end
      end else begin
        if(when_DCache_l237_1) begin
          if(cache_hit_1) begin
            if(_zz_12) begin
              ways_1_metas_0_mru <= 1'b1;
            end
            if(_zz_13) begin
              ways_1_metas_1_mru <= 1'b1;
            end
            if(_zz_14) begin
              ways_1_metas_2_mru <= 1'b1;
            end
            if(_zz_15) begin
              ways_1_metas_3_mru <= 1'b1;
            end
          end else begin
            if(_zz_12) begin
              ways_1_metas_0_mru <= 1'b0;
            end
            if(_zz_13) begin
              ways_1_metas_1_mru <= 1'b0;
            end
            if(_zz_14) begin
              ways_1_metas_2_mru <= 1'b0;
            end
            if(_zz_15) begin
              ways_1_metas_3_mru <= 1'b0;
            end
          end
        end else begin
          if(when_DCache_l244_1) begin
            if(_zz_12) begin
              ways_1_metas_0_mru <= 1'b1;
            end
            if(_zz_13) begin
              ways_1_metas_1_mru <= 1'b1;
            end
            if(_zz_14) begin
              ways_1_metas_2_mru <= 1'b1;
            end
            if(_zz_15) begin
              ways_1_metas_3_mru <= 1'b1;
            end
          end else begin
            if(when_DCache_l247_1) begin
              if(_zz_12) begin
                ways_1_metas_0_vld <= 1'b1;
              end
              if(_zz_13) begin
                ways_1_metas_1_vld <= 1'b1;
              end
              if(_zz_14) begin
                ways_1_metas_2_vld <= 1'b1;
              end
              if(_zz_15) begin
                ways_1_metas_3_vld <= 1'b1;
              end
            end
          end
        end
      end
      if(when_DCache_l252_1) begin
        if(_zz_12) begin
          ways_1_metas_0_tag <= cpu_tag;
        end
        if(_zz_13) begin
          ways_1_metas_1_tag <= cpu_tag;
        end
        if(_zz_14) begin
          ways_1_metas_2_tag <= cpu_tag;
        end
        if(_zz_15) begin
          ways_1_metas_3_tag <= cpu_tag;
        end
      end
      if(flush_busy) begin
        if(_zz_27) begin
          ways_2_metas_0_mru <= 1'b0;
        end
        if(_zz_28) begin
          ways_2_metas_1_mru <= 1'b0;
        end
        if(_zz_29) begin
          ways_2_metas_2_mru <= 1'b0;
        end
        if(_zz_30) begin
          ways_2_metas_3_mru <= 1'b0;
        end
        if(_zz_27) begin
          ways_2_metas_0_vld <= 1'b0;
        end
        if(_zz_28) begin
          ways_2_metas_1_vld <= 1'b0;
        end
        if(_zz_29) begin
          ways_2_metas_2_vld <= 1'b0;
        end
        if(_zz_30) begin
          ways_2_metas_3_vld <= 1'b0;
        end
      end else begin
        if(when_DCache_l237_2) begin
          if(cache_hit_2) begin
            if(_zz_22) begin
              ways_2_metas_0_mru <= 1'b1;
            end
            if(_zz_23) begin
              ways_2_metas_1_mru <= 1'b1;
            end
            if(_zz_24) begin
              ways_2_metas_2_mru <= 1'b1;
            end
            if(_zz_25) begin
              ways_2_metas_3_mru <= 1'b1;
            end
          end else begin
            if(_zz_22) begin
              ways_2_metas_0_mru <= 1'b0;
            end
            if(_zz_23) begin
              ways_2_metas_1_mru <= 1'b0;
            end
            if(_zz_24) begin
              ways_2_metas_2_mru <= 1'b0;
            end
            if(_zz_25) begin
              ways_2_metas_3_mru <= 1'b0;
            end
          end
        end else begin
          if(when_DCache_l244_2) begin
            if(_zz_22) begin
              ways_2_metas_0_mru <= 1'b1;
            end
            if(_zz_23) begin
              ways_2_metas_1_mru <= 1'b1;
            end
            if(_zz_24) begin
              ways_2_metas_2_mru <= 1'b1;
            end
            if(_zz_25) begin
              ways_2_metas_3_mru <= 1'b1;
            end
          end else begin
            if(when_DCache_l247_2) begin
              if(_zz_22) begin
                ways_2_metas_0_vld <= 1'b1;
              end
              if(_zz_23) begin
                ways_2_metas_1_vld <= 1'b1;
              end
              if(_zz_24) begin
                ways_2_metas_2_vld <= 1'b1;
              end
              if(_zz_25) begin
                ways_2_metas_3_vld <= 1'b1;
              end
            end
          end
        end
      end
      if(when_DCache_l252_2) begin
        if(_zz_22) begin
          ways_2_metas_0_tag <= cpu_tag;
        end
        if(_zz_23) begin
          ways_2_metas_1_tag <= cpu_tag;
        end
        if(_zz_24) begin
          ways_2_metas_2_tag <= cpu_tag;
        end
        if(_zz_25) begin
          ways_2_metas_3_tag <= cpu_tag;
        end
      end
      if(flush_busy) begin
        if(_zz_37) begin
          ways_3_metas_0_mru <= 1'b0;
        end
        if(_zz_38) begin
          ways_3_metas_1_mru <= 1'b0;
        end
        if(_zz_39) begin
          ways_3_metas_2_mru <= 1'b0;
        end
        if(_zz_40) begin
          ways_3_metas_3_mru <= 1'b0;
        end
        if(_zz_37) begin
          ways_3_metas_0_vld <= 1'b0;
        end
        if(_zz_38) begin
          ways_3_metas_1_vld <= 1'b0;
        end
        if(_zz_39) begin
          ways_3_metas_2_vld <= 1'b0;
        end
        if(_zz_40) begin
          ways_3_metas_3_vld <= 1'b0;
        end
      end else begin
        if(when_DCache_l237_3) begin
          if(cache_hit_3) begin
            if(_zz_32) begin
              ways_3_metas_0_mru <= 1'b1;
            end
            if(_zz_33) begin
              ways_3_metas_1_mru <= 1'b1;
            end
            if(_zz_34) begin
              ways_3_metas_2_mru <= 1'b1;
            end
            if(_zz_35) begin
              ways_3_metas_3_mru <= 1'b1;
            end
          end else begin
            if(_zz_32) begin
              ways_3_metas_0_mru <= 1'b0;
            end
            if(_zz_33) begin
              ways_3_metas_1_mru <= 1'b0;
            end
            if(_zz_34) begin
              ways_3_metas_2_mru <= 1'b0;
            end
            if(_zz_35) begin
              ways_3_metas_3_mru <= 1'b0;
            end
          end
        end else begin
          if(when_DCache_l244_3) begin
            if(_zz_32) begin
              ways_3_metas_0_mru <= 1'b1;
            end
            if(_zz_33) begin
              ways_3_metas_1_mru <= 1'b1;
            end
            if(_zz_34) begin
              ways_3_metas_2_mru <= 1'b1;
            end
            if(_zz_35) begin
              ways_3_metas_3_mru <= 1'b1;
            end
          end else begin
            if(when_DCache_l247_3) begin
              if(_zz_32) begin
                ways_3_metas_0_vld <= 1'b1;
              end
              if(_zz_33) begin
                ways_3_metas_1_vld <= 1'b1;
              end
              if(_zz_34) begin
                ways_3_metas_2_vld <= 1'b1;
              end
              if(_zz_35) begin
                ways_3_metas_3_vld <= 1'b1;
              end
            end
          end
        end
      end
      if(when_DCache_l252_3) begin
        if(_zz_32) begin
          ways_3_metas_0_tag <= cpu_tag;
        end
        if(_zz_33) begin
          ways_3_metas_1_tag <= cpu_tag;
        end
        if(_zz_34) begin
          ways_3_metas_2_tag <= cpu_tag;
        end
        if(_zz_35) begin
          ways_3_metas_3_tag <= cpu_tag;
        end
      end
      if(when_DCache_l258) begin
        cpu_cmd_ready_1 <= 1'b0;
      end else begin
        if(when_DCache_l261) begin
          cpu_cmd_ready_1 <= 1'b1;
        end
      end
    end
  end

  always @(posedge io_axiClk) begin
    bypass_rsp_valid_d1 <= cpu_bypass_rsp_valid;
    bypass_rsp_data_d1 <= cpu_bypass_rsp_payload_data;
    if(is_miss) begin
      evict_id_miss <= evict_id;
    end
    next_level_rdone <= (next_level_rvalid && (next_level_data_cnt_value == 3'b111));
    next_level_wdone <= ((next_level_rsp_valid && (! next_level_rsp_payload_rvalid)) && (next_level_rsp_payload_bresp == 2'b00));
  end


endmodule

module SramBanks (
  input               sram_0_ports_cmd_valid,
  input      [3:0]    sram_0_ports_cmd_payload_addr,
  input      [15:0]   sram_0_ports_cmd_payload_wen,
  input      [511:0]  sram_0_ports_cmd_payload_wdata,
  input      [63:0]   sram_0_ports_cmd_payload_wstrb,
  output              sram_0_ports_rsp_valid,
  output reg [511:0]  sram_0_ports_rsp_payload_data,
  input               sram_1_ports_cmd_valid,
  input      [3:0]    sram_1_ports_cmd_payload_addr,
  input      [15:0]   sram_1_ports_cmd_payload_wen,
  input      [511:0]  sram_1_ports_cmd_payload_wdata,
  input      [63:0]   sram_1_ports_cmd_payload_wstrb,
  output              sram_1_ports_rsp_valid,
  output reg [511:0]  sram_1_ports_rsp_payload_data,
  input               sram_2_ports_cmd_valid,
  input      [3:0]    sram_2_ports_cmd_payload_addr,
  input      [15:0]   sram_2_ports_cmd_payload_wen,
  input      [511:0]  sram_2_ports_cmd_payload_wdata,
  input      [63:0]   sram_2_ports_cmd_payload_wstrb,
  output              sram_2_ports_rsp_valid,
  output reg [511:0]  sram_2_ports_rsp_payload_data,
  input               sram_3_ports_cmd_valid,
  input      [3:0]    sram_3_ports_cmd_payload_addr,
  input      [15:0]   sram_3_ports_cmd_payload_wen,
  input      [511:0]  sram_3_ports_cmd_payload_wdata,
  input      [63:0]   sram_3_ports_cmd_payload_wstrb,
  output              sram_3_ports_rsp_valid,
  output reg [511:0]  sram_3_ports_rsp_payload_data,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  reg        [31:0]   _zz_sram_0_banks_0_bank_port1;
  reg        [31:0]   _zz_sram_0_banks_1_bank_port1;
  reg        [31:0]   _zz_sram_0_banks_2_bank_port1;
  reg        [31:0]   _zz_sram_0_banks_3_bank_port1;
  reg        [31:0]   _zz_sram_0_banks_4_bank_port1;
  reg        [31:0]   _zz_sram_0_banks_5_bank_port1;
  reg        [31:0]   _zz_sram_0_banks_6_bank_port1;
  reg        [31:0]   _zz_sram_0_banks_7_bank_port1;
  reg        [31:0]   _zz_sram_0_banks_8_bank_port1;
  reg        [31:0]   _zz_sram_0_banks_9_bank_port1;
  reg        [31:0]   _zz_sram_0_banks_10_bank_port1;
  reg        [31:0]   _zz_sram_0_banks_11_bank_port1;
  reg        [31:0]   _zz_sram_0_banks_12_bank_port1;
  reg        [31:0]   _zz_sram_0_banks_13_bank_port1;
  reg        [31:0]   _zz_sram_0_banks_14_bank_port1;
  reg        [31:0]   _zz_sram_0_banks_15_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_0_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_1_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_2_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_3_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_4_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_5_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_6_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_7_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_8_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_9_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_10_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_11_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_12_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_13_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_14_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_15_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_0_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_1_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_2_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_3_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_4_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_5_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_6_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_7_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_8_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_9_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_10_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_11_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_12_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_13_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_14_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_15_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_0_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_1_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_2_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_3_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_4_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_5_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_6_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_7_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_8_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_9_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_10_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_11_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_12_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_13_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_14_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_15_bank_port1;
  wire       [31:0]   _zz_sram_0_banks_0_bank_port;
  wire       [3:0]    _zz_sram_0_banks_0_bank_port_1;
  wire                _zz_sram_0_banks_0_bank_port_2;
  wire       [31:0]   _zz_sram_0_banks_1_bank_port;
  wire       [3:0]    _zz_sram_0_banks_1_bank_port_1;
  wire                _zz_sram_0_banks_1_bank_port_2;
  wire       [31:0]   _zz_sram_0_banks_2_bank_port;
  wire       [3:0]    _zz_sram_0_banks_2_bank_port_1;
  wire                _zz_sram_0_banks_2_bank_port_2;
  wire       [31:0]   _zz_sram_0_banks_3_bank_port;
  wire       [3:0]    _zz_sram_0_banks_3_bank_port_1;
  wire                _zz_sram_0_banks_3_bank_port_2;
  wire       [31:0]   _zz_sram_0_banks_4_bank_port;
  wire       [3:0]    _zz_sram_0_banks_4_bank_port_1;
  wire                _zz_sram_0_banks_4_bank_port_2;
  wire       [31:0]   _zz_sram_0_banks_5_bank_port;
  wire       [3:0]    _zz_sram_0_banks_5_bank_port_1;
  wire                _zz_sram_0_banks_5_bank_port_2;
  wire       [31:0]   _zz_sram_0_banks_6_bank_port;
  wire       [3:0]    _zz_sram_0_banks_6_bank_port_1;
  wire                _zz_sram_0_banks_6_bank_port_2;
  wire       [31:0]   _zz_sram_0_banks_7_bank_port;
  wire       [3:0]    _zz_sram_0_banks_7_bank_port_1;
  wire                _zz_sram_0_banks_7_bank_port_2;
  wire       [31:0]   _zz_sram_0_banks_8_bank_port;
  wire       [3:0]    _zz_sram_0_banks_8_bank_port_1;
  wire                _zz_sram_0_banks_8_bank_port_2;
  wire       [31:0]   _zz_sram_0_banks_9_bank_port;
  wire       [3:0]    _zz_sram_0_banks_9_bank_port_1;
  wire                _zz_sram_0_banks_9_bank_port_2;
  wire       [31:0]   _zz_sram_0_banks_10_bank_port;
  wire       [3:0]    _zz_sram_0_banks_10_bank_port_1;
  wire                _zz_sram_0_banks_10_bank_port_2;
  wire       [31:0]   _zz_sram_0_banks_11_bank_port;
  wire       [3:0]    _zz_sram_0_banks_11_bank_port_1;
  wire                _zz_sram_0_banks_11_bank_port_2;
  wire       [31:0]   _zz_sram_0_banks_12_bank_port;
  wire       [3:0]    _zz_sram_0_banks_12_bank_port_1;
  wire                _zz_sram_0_banks_12_bank_port_2;
  wire       [31:0]   _zz_sram_0_banks_13_bank_port;
  wire       [3:0]    _zz_sram_0_banks_13_bank_port_1;
  wire                _zz_sram_0_banks_13_bank_port_2;
  wire       [31:0]   _zz_sram_0_banks_14_bank_port;
  wire       [3:0]    _zz_sram_0_banks_14_bank_port_1;
  wire                _zz_sram_0_banks_14_bank_port_2;
  wire       [31:0]   _zz_sram_0_banks_15_bank_port;
  wire       [3:0]    _zz_sram_0_banks_15_bank_port_1;
  wire                _zz_sram_0_banks_15_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_0_bank_port;
  wire       [3:0]    _zz_sram_1_banks_0_bank_port_1;
  wire                _zz_sram_1_banks_0_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_1_bank_port;
  wire       [3:0]    _zz_sram_1_banks_1_bank_port_1;
  wire                _zz_sram_1_banks_1_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_2_bank_port;
  wire       [3:0]    _zz_sram_1_banks_2_bank_port_1;
  wire                _zz_sram_1_banks_2_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_3_bank_port;
  wire       [3:0]    _zz_sram_1_banks_3_bank_port_1;
  wire                _zz_sram_1_banks_3_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_4_bank_port;
  wire       [3:0]    _zz_sram_1_banks_4_bank_port_1;
  wire                _zz_sram_1_banks_4_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_5_bank_port;
  wire       [3:0]    _zz_sram_1_banks_5_bank_port_1;
  wire                _zz_sram_1_banks_5_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_6_bank_port;
  wire       [3:0]    _zz_sram_1_banks_6_bank_port_1;
  wire                _zz_sram_1_banks_6_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_7_bank_port;
  wire       [3:0]    _zz_sram_1_banks_7_bank_port_1;
  wire                _zz_sram_1_banks_7_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_8_bank_port;
  wire       [3:0]    _zz_sram_1_banks_8_bank_port_1;
  wire                _zz_sram_1_banks_8_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_9_bank_port;
  wire       [3:0]    _zz_sram_1_banks_9_bank_port_1;
  wire                _zz_sram_1_banks_9_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_10_bank_port;
  wire       [3:0]    _zz_sram_1_banks_10_bank_port_1;
  wire                _zz_sram_1_banks_10_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_11_bank_port;
  wire       [3:0]    _zz_sram_1_banks_11_bank_port_1;
  wire                _zz_sram_1_banks_11_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_12_bank_port;
  wire       [3:0]    _zz_sram_1_banks_12_bank_port_1;
  wire                _zz_sram_1_banks_12_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_13_bank_port;
  wire       [3:0]    _zz_sram_1_banks_13_bank_port_1;
  wire                _zz_sram_1_banks_13_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_14_bank_port;
  wire       [3:0]    _zz_sram_1_banks_14_bank_port_1;
  wire                _zz_sram_1_banks_14_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_15_bank_port;
  wire       [3:0]    _zz_sram_1_banks_15_bank_port_1;
  wire                _zz_sram_1_banks_15_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_0_bank_port;
  wire       [3:0]    _zz_sram_2_banks_0_bank_port_1;
  wire                _zz_sram_2_banks_0_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_1_bank_port;
  wire       [3:0]    _zz_sram_2_banks_1_bank_port_1;
  wire                _zz_sram_2_banks_1_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_2_bank_port;
  wire       [3:0]    _zz_sram_2_banks_2_bank_port_1;
  wire                _zz_sram_2_banks_2_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_3_bank_port;
  wire       [3:0]    _zz_sram_2_banks_3_bank_port_1;
  wire                _zz_sram_2_banks_3_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_4_bank_port;
  wire       [3:0]    _zz_sram_2_banks_4_bank_port_1;
  wire                _zz_sram_2_banks_4_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_5_bank_port;
  wire       [3:0]    _zz_sram_2_banks_5_bank_port_1;
  wire                _zz_sram_2_banks_5_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_6_bank_port;
  wire       [3:0]    _zz_sram_2_banks_6_bank_port_1;
  wire                _zz_sram_2_banks_6_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_7_bank_port;
  wire       [3:0]    _zz_sram_2_banks_7_bank_port_1;
  wire                _zz_sram_2_banks_7_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_8_bank_port;
  wire       [3:0]    _zz_sram_2_banks_8_bank_port_1;
  wire                _zz_sram_2_banks_8_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_9_bank_port;
  wire       [3:0]    _zz_sram_2_banks_9_bank_port_1;
  wire                _zz_sram_2_banks_9_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_10_bank_port;
  wire       [3:0]    _zz_sram_2_banks_10_bank_port_1;
  wire                _zz_sram_2_banks_10_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_11_bank_port;
  wire       [3:0]    _zz_sram_2_banks_11_bank_port_1;
  wire                _zz_sram_2_banks_11_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_12_bank_port;
  wire       [3:0]    _zz_sram_2_banks_12_bank_port_1;
  wire                _zz_sram_2_banks_12_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_13_bank_port;
  wire       [3:0]    _zz_sram_2_banks_13_bank_port_1;
  wire                _zz_sram_2_banks_13_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_14_bank_port;
  wire       [3:0]    _zz_sram_2_banks_14_bank_port_1;
  wire                _zz_sram_2_banks_14_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_15_bank_port;
  wire       [3:0]    _zz_sram_2_banks_15_bank_port_1;
  wire                _zz_sram_2_banks_15_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_0_bank_port;
  wire       [3:0]    _zz_sram_3_banks_0_bank_port_1;
  wire                _zz_sram_3_banks_0_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_1_bank_port;
  wire       [3:0]    _zz_sram_3_banks_1_bank_port_1;
  wire                _zz_sram_3_banks_1_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_2_bank_port;
  wire       [3:0]    _zz_sram_3_banks_2_bank_port_1;
  wire                _zz_sram_3_banks_2_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_3_bank_port;
  wire       [3:0]    _zz_sram_3_banks_3_bank_port_1;
  wire                _zz_sram_3_banks_3_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_4_bank_port;
  wire       [3:0]    _zz_sram_3_banks_4_bank_port_1;
  wire                _zz_sram_3_banks_4_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_5_bank_port;
  wire       [3:0]    _zz_sram_3_banks_5_bank_port_1;
  wire                _zz_sram_3_banks_5_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_6_bank_port;
  wire       [3:0]    _zz_sram_3_banks_6_bank_port_1;
  wire                _zz_sram_3_banks_6_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_7_bank_port;
  wire       [3:0]    _zz_sram_3_banks_7_bank_port_1;
  wire                _zz_sram_3_banks_7_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_8_bank_port;
  wire       [3:0]    _zz_sram_3_banks_8_bank_port_1;
  wire                _zz_sram_3_banks_8_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_9_bank_port;
  wire       [3:0]    _zz_sram_3_banks_9_bank_port_1;
  wire                _zz_sram_3_banks_9_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_10_bank_port;
  wire       [3:0]    _zz_sram_3_banks_10_bank_port_1;
  wire                _zz_sram_3_banks_10_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_11_bank_port;
  wire       [3:0]    _zz_sram_3_banks_11_bank_port_1;
  wire                _zz_sram_3_banks_11_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_12_bank_port;
  wire       [3:0]    _zz_sram_3_banks_12_bank_port_1;
  wire                _zz_sram_3_banks_12_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_13_bank_port;
  wire       [3:0]    _zz_sram_3_banks_13_bank_port_1;
  wire                _zz_sram_3_banks_13_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_14_bank_port;
  wire       [3:0]    _zz_sram_3_banks_14_bank_port_1;
  wire                _zz_sram_3_banks_14_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_15_bank_port;
  wire       [3:0]    _zz_sram_3_banks_15_bank_port_1;
  wire                _zz_sram_3_banks_15_bank_port_2;
  reg                 _zz_sram_0_ports_rsp_valid;
  wire                when_SramBanks_l66;
  reg                 _zz_sram_1_ports_rsp_valid;
  wire                when_SramBanks_l66_1;
  reg                 _zz_sram_2_ports_rsp_valid;
  wire                when_SramBanks_l66_2;
  reg                 _zz_sram_3_ports_rsp_valid;
  wire                when_SramBanks_l66_3;
  reg [7:0] sram_0_banks_0_bank_symbol0 [0:15];
  reg [7:0] sram_0_banks_0_bank_symbol1 [0:15];
  reg [7:0] sram_0_banks_0_bank_symbol2 [0:15];
  reg [7:0] sram_0_banks_0_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_0_banks_0_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_0_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_0_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_0_banksymbol_read_3;
  reg [7:0] sram_0_banks_1_bank_symbol0 [0:15];
  reg [7:0] sram_0_banks_1_bank_symbol1 [0:15];
  reg [7:0] sram_0_banks_1_bank_symbol2 [0:15];
  reg [7:0] sram_0_banks_1_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_0_banks_1_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_1_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_1_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_1_banksymbol_read_3;
  reg [7:0] sram_0_banks_2_bank_symbol0 [0:15];
  reg [7:0] sram_0_banks_2_bank_symbol1 [0:15];
  reg [7:0] sram_0_banks_2_bank_symbol2 [0:15];
  reg [7:0] sram_0_banks_2_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_0_banks_2_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_2_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_2_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_2_banksymbol_read_3;
  reg [7:0] sram_0_banks_3_bank_symbol0 [0:15];
  reg [7:0] sram_0_banks_3_bank_symbol1 [0:15];
  reg [7:0] sram_0_banks_3_bank_symbol2 [0:15];
  reg [7:0] sram_0_banks_3_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_0_banks_3_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_3_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_3_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_3_banksymbol_read_3;
  reg [7:0] sram_0_banks_4_bank_symbol0 [0:15];
  reg [7:0] sram_0_banks_4_bank_symbol1 [0:15];
  reg [7:0] sram_0_banks_4_bank_symbol2 [0:15];
  reg [7:0] sram_0_banks_4_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_0_banks_4_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_4_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_4_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_4_banksymbol_read_3;
  reg [7:0] sram_0_banks_5_bank_symbol0 [0:15];
  reg [7:0] sram_0_banks_5_bank_symbol1 [0:15];
  reg [7:0] sram_0_banks_5_bank_symbol2 [0:15];
  reg [7:0] sram_0_banks_5_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_0_banks_5_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_5_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_5_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_5_banksymbol_read_3;
  reg [7:0] sram_0_banks_6_bank_symbol0 [0:15];
  reg [7:0] sram_0_banks_6_bank_symbol1 [0:15];
  reg [7:0] sram_0_banks_6_bank_symbol2 [0:15];
  reg [7:0] sram_0_banks_6_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_0_banks_6_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_6_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_6_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_6_banksymbol_read_3;
  reg [7:0] sram_0_banks_7_bank_symbol0 [0:15];
  reg [7:0] sram_0_banks_7_bank_symbol1 [0:15];
  reg [7:0] sram_0_banks_7_bank_symbol2 [0:15];
  reg [7:0] sram_0_banks_7_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_0_banks_7_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_7_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_7_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_7_banksymbol_read_3;
  reg [7:0] sram_0_banks_8_bank_symbol0 [0:15];
  reg [7:0] sram_0_banks_8_bank_symbol1 [0:15];
  reg [7:0] sram_0_banks_8_bank_symbol2 [0:15];
  reg [7:0] sram_0_banks_8_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_0_banks_8_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_8_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_8_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_8_banksymbol_read_3;
  reg [7:0] sram_0_banks_9_bank_symbol0 [0:15];
  reg [7:0] sram_0_banks_9_bank_symbol1 [0:15];
  reg [7:0] sram_0_banks_9_bank_symbol2 [0:15];
  reg [7:0] sram_0_banks_9_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_0_banks_9_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_9_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_9_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_9_banksymbol_read_3;
  reg [7:0] sram_0_banks_10_bank_symbol0 [0:15];
  reg [7:0] sram_0_banks_10_bank_symbol1 [0:15];
  reg [7:0] sram_0_banks_10_bank_symbol2 [0:15];
  reg [7:0] sram_0_banks_10_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_0_banks_10_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_10_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_10_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_10_banksymbol_read_3;
  reg [7:0] sram_0_banks_11_bank_symbol0 [0:15];
  reg [7:0] sram_0_banks_11_bank_symbol1 [0:15];
  reg [7:0] sram_0_banks_11_bank_symbol2 [0:15];
  reg [7:0] sram_0_banks_11_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_0_banks_11_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_11_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_11_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_11_banksymbol_read_3;
  reg [7:0] sram_0_banks_12_bank_symbol0 [0:15];
  reg [7:0] sram_0_banks_12_bank_symbol1 [0:15];
  reg [7:0] sram_0_banks_12_bank_symbol2 [0:15];
  reg [7:0] sram_0_banks_12_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_0_banks_12_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_12_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_12_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_12_banksymbol_read_3;
  reg [7:0] sram_0_banks_13_bank_symbol0 [0:15];
  reg [7:0] sram_0_banks_13_bank_symbol1 [0:15];
  reg [7:0] sram_0_banks_13_bank_symbol2 [0:15];
  reg [7:0] sram_0_banks_13_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_0_banks_13_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_13_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_13_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_13_banksymbol_read_3;
  reg [7:0] sram_0_banks_14_bank_symbol0 [0:15];
  reg [7:0] sram_0_banks_14_bank_symbol1 [0:15];
  reg [7:0] sram_0_banks_14_bank_symbol2 [0:15];
  reg [7:0] sram_0_banks_14_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_0_banks_14_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_14_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_14_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_14_banksymbol_read_3;
  reg [7:0] sram_0_banks_15_bank_symbol0 [0:15];
  reg [7:0] sram_0_banks_15_bank_symbol1 [0:15];
  reg [7:0] sram_0_banks_15_bank_symbol2 [0:15];
  reg [7:0] sram_0_banks_15_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_0_banks_15_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_15_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_15_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_15_banksymbol_read_3;
  reg [7:0] sram_1_banks_0_bank_symbol0 [0:15];
  reg [7:0] sram_1_banks_0_bank_symbol1 [0:15];
  reg [7:0] sram_1_banks_0_bank_symbol2 [0:15];
  reg [7:0] sram_1_banks_0_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_1_banks_0_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_0_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_0_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_0_banksymbol_read_3;
  reg [7:0] sram_1_banks_1_bank_symbol0 [0:15];
  reg [7:0] sram_1_banks_1_bank_symbol1 [0:15];
  reg [7:0] sram_1_banks_1_bank_symbol2 [0:15];
  reg [7:0] sram_1_banks_1_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_1_banks_1_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_1_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_1_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_1_banksymbol_read_3;
  reg [7:0] sram_1_banks_2_bank_symbol0 [0:15];
  reg [7:0] sram_1_banks_2_bank_symbol1 [0:15];
  reg [7:0] sram_1_banks_2_bank_symbol2 [0:15];
  reg [7:0] sram_1_banks_2_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_1_banks_2_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_2_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_2_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_2_banksymbol_read_3;
  reg [7:0] sram_1_banks_3_bank_symbol0 [0:15];
  reg [7:0] sram_1_banks_3_bank_symbol1 [0:15];
  reg [7:0] sram_1_banks_3_bank_symbol2 [0:15];
  reg [7:0] sram_1_banks_3_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_1_banks_3_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_3_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_3_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_3_banksymbol_read_3;
  reg [7:0] sram_1_banks_4_bank_symbol0 [0:15];
  reg [7:0] sram_1_banks_4_bank_symbol1 [0:15];
  reg [7:0] sram_1_banks_4_bank_symbol2 [0:15];
  reg [7:0] sram_1_banks_4_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_1_banks_4_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_4_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_4_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_4_banksymbol_read_3;
  reg [7:0] sram_1_banks_5_bank_symbol0 [0:15];
  reg [7:0] sram_1_banks_5_bank_symbol1 [0:15];
  reg [7:0] sram_1_banks_5_bank_symbol2 [0:15];
  reg [7:0] sram_1_banks_5_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_1_banks_5_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_5_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_5_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_5_banksymbol_read_3;
  reg [7:0] sram_1_banks_6_bank_symbol0 [0:15];
  reg [7:0] sram_1_banks_6_bank_symbol1 [0:15];
  reg [7:0] sram_1_banks_6_bank_symbol2 [0:15];
  reg [7:0] sram_1_banks_6_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_1_banks_6_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_6_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_6_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_6_banksymbol_read_3;
  reg [7:0] sram_1_banks_7_bank_symbol0 [0:15];
  reg [7:0] sram_1_banks_7_bank_symbol1 [0:15];
  reg [7:0] sram_1_banks_7_bank_symbol2 [0:15];
  reg [7:0] sram_1_banks_7_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_1_banks_7_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_7_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_7_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_7_banksymbol_read_3;
  reg [7:0] sram_1_banks_8_bank_symbol0 [0:15];
  reg [7:0] sram_1_banks_8_bank_symbol1 [0:15];
  reg [7:0] sram_1_banks_8_bank_symbol2 [0:15];
  reg [7:0] sram_1_banks_8_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_1_banks_8_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_8_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_8_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_8_banksymbol_read_3;
  reg [7:0] sram_1_banks_9_bank_symbol0 [0:15];
  reg [7:0] sram_1_banks_9_bank_symbol1 [0:15];
  reg [7:0] sram_1_banks_9_bank_symbol2 [0:15];
  reg [7:0] sram_1_banks_9_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_1_banks_9_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_9_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_9_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_9_banksymbol_read_3;
  reg [7:0] sram_1_banks_10_bank_symbol0 [0:15];
  reg [7:0] sram_1_banks_10_bank_symbol1 [0:15];
  reg [7:0] sram_1_banks_10_bank_symbol2 [0:15];
  reg [7:0] sram_1_banks_10_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_1_banks_10_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_10_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_10_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_10_banksymbol_read_3;
  reg [7:0] sram_1_banks_11_bank_symbol0 [0:15];
  reg [7:0] sram_1_banks_11_bank_symbol1 [0:15];
  reg [7:0] sram_1_banks_11_bank_symbol2 [0:15];
  reg [7:0] sram_1_banks_11_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_1_banks_11_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_11_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_11_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_11_banksymbol_read_3;
  reg [7:0] sram_1_banks_12_bank_symbol0 [0:15];
  reg [7:0] sram_1_banks_12_bank_symbol1 [0:15];
  reg [7:0] sram_1_banks_12_bank_symbol2 [0:15];
  reg [7:0] sram_1_banks_12_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_1_banks_12_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_12_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_12_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_12_banksymbol_read_3;
  reg [7:0] sram_1_banks_13_bank_symbol0 [0:15];
  reg [7:0] sram_1_banks_13_bank_symbol1 [0:15];
  reg [7:0] sram_1_banks_13_bank_symbol2 [0:15];
  reg [7:0] sram_1_banks_13_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_1_banks_13_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_13_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_13_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_13_banksymbol_read_3;
  reg [7:0] sram_1_banks_14_bank_symbol0 [0:15];
  reg [7:0] sram_1_banks_14_bank_symbol1 [0:15];
  reg [7:0] sram_1_banks_14_bank_symbol2 [0:15];
  reg [7:0] sram_1_banks_14_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_1_banks_14_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_14_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_14_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_14_banksymbol_read_3;
  reg [7:0] sram_1_banks_15_bank_symbol0 [0:15];
  reg [7:0] sram_1_banks_15_bank_symbol1 [0:15];
  reg [7:0] sram_1_banks_15_bank_symbol2 [0:15];
  reg [7:0] sram_1_banks_15_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_1_banks_15_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_15_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_15_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_15_banksymbol_read_3;
  reg [7:0] sram_2_banks_0_bank_symbol0 [0:15];
  reg [7:0] sram_2_banks_0_bank_symbol1 [0:15];
  reg [7:0] sram_2_banks_0_bank_symbol2 [0:15];
  reg [7:0] sram_2_banks_0_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_2_banks_0_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_0_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_0_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_0_banksymbol_read_3;
  reg [7:0] sram_2_banks_1_bank_symbol0 [0:15];
  reg [7:0] sram_2_banks_1_bank_symbol1 [0:15];
  reg [7:0] sram_2_banks_1_bank_symbol2 [0:15];
  reg [7:0] sram_2_banks_1_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_2_banks_1_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_1_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_1_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_1_banksymbol_read_3;
  reg [7:0] sram_2_banks_2_bank_symbol0 [0:15];
  reg [7:0] sram_2_banks_2_bank_symbol1 [0:15];
  reg [7:0] sram_2_banks_2_bank_symbol2 [0:15];
  reg [7:0] sram_2_banks_2_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_2_banks_2_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_2_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_2_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_2_banksymbol_read_3;
  reg [7:0] sram_2_banks_3_bank_symbol0 [0:15];
  reg [7:0] sram_2_banks_3_bank_symbol1 [0:15];
  reg [7:0] sram_2_banks_3_bank_symbol2 [0:15];
  reg [7:0] sram_2_banks_3_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_2_banks_3_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_3_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_3_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_3_banksymbol_read_3;
  reg [7:0] sram_2_banks_4_bank_symbol0 [0:15];
  reg [7:0] sram_2_banks_4_bank_symbol1 [0:15];
  reg [7:0] sram_2_banks_4_bank_symbol2 [0:15];
  reg [7:0] sram_2_banks_4_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_2_banks_4_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_4_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_4_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_4_banksymbol_read_3;
  reg [7:0] sram_2_banks_5_bank_symbol0 [0:15];
  reg [7:0] sram_2_banks_5_bank_symbol1 [0:15];
  reg [7:0] sram_2_banks_5_bank_symbol2 [0:15];
  reg [7:0] sram_2_banks_5_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_2_banks_5_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_5_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_5_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_5_banksymbol_read_3;
  reg [7:0] sram_2_banks_6_bank_symbol0 [0:15];
  reg [7:0] sram_2_banks_6_bank_symbol1 [0:15];
  reg [7:0] sram_2_banks_6_bank_symbol2 [0:15];
  reg [7:0] sram_2_banks_6_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_2_banks_6_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_6_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_6_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_6_banksymbol_read_3;
  reg [7:0] sram_2_banks_7_bank_symbol0 [0:15];
  reg [7:0] sram_2_banks_7_bank_symbol1 [0:15];
  reg [7:0] sram_2_banks_7_bank_symbol2 [0:15];
  reg [7:0] sram_2_banks_7_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_2_banks_7_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_7_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_7_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_7_banksymbol_read_3;
  reg [7:0] sram_2_banks_8_bank_symbol0 [0:15];
  reg [7:0] sram_2_banks_8_bank_symbol1 [0:15];
  reg [7:0] sram_2_banks_8_bank_symbol2 [0:15];
  reg [7:0] sram_2_banks_8_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_2_banks_8_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_8_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_8_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_8_banksymbol_read_3;
  reg [7:0] sram_2_banks_9_bank_symbol0 [0:15];
  reg [7:0] sram_2_banks_9_bank_symbol1 [0:15];
  reg [7:0] sram_2_banks_9_bank_symbol2 [0:15];
  reg [7:0] sram_2_banks_9_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_2_banks_9_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_9_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_9_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_9_banksymbol_read_3;
  reg [7:0] sram_2_banks_10_bank_symbol0 [0:15];
  reg [7:0] sram_2_banks_10_bank_symbol1 [0:15];
  reg [7:0] sram_2_banks_10_bank_symbol2 [0:15];
  reg [7:0] sram_2_banks_10_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_2_banks_10_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_10_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_10_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_10_banksymbol_read_3;
  reg [7:0] sram_2_banks_11_bank_symbol0 [0:15];
  reg [7:0] sram_2_banks_11_bank_symbol1 [0:15];
  reg [7:0] sram_2_banks_11_bank_symbol2 [0:15];
  reg [7:0] sram_2_banks_11_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_2_banks_11_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_11_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_11_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_11_banksymbol_read_3;
  reg [7:0] sram_2_banks_12_bank_symbol0 [0:15];
  reg [7:0] sram_2_banks_12_bank_symbol1 [0:15];
  reg [7:0] sram_2_banks_12_bank_symbol2 [0:15];
  reg [7:0] sram_2_banks_12_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_2_banks_12_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_12_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_12_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_12_banksymbol_read_3;
  reg [7:0] sram_2_banks_13_bank_symbol0 [0:15];
  reg [7:0] sram_2_banks_13_bank_symbol1 [0:15];
  reg [7:0] sram_2_banks_13_bank_symbol2 [0:15];
  reg [7:0] sram_2_banks_13_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_2_banks_13_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_13_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_13_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_13_banksymbol_read_3;
  reg [7:0] sram_2_banks_14_bank_symbol0 [0:15];
  reg [7:0] sram_2_banks_14_bank_symbol1 [0:15];
  reg [7:0] sram_2_banks_14_bank_symbol2 [0:15];
  reg [7:0] sram_2_banks_14_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_2_banks_14_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_14_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_14_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_14_banksymbol_read_3;
  reg [7:0] sram_2_banks_15_bank_symbol0 [0:15];
  reg [7:0] sram_2_banks_15_bank_symbol1 [0:15];
  reg [7:0] sram_2_banks_15_bank_symbol2 [0:15];
  reg [7:0] sram_2_banks_15_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_2_banks_15_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_15_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_15_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_15_banksymbol_read_3;
  reg [7:0] sram_3_banks_0_bank_symbol0 [0:15];
  reg [7:0] sram_3_banks_0_bank_symbol1 [0:15];
  reg [7:0] sram_3_banks_0_bank_symbol2 [0:15];
  reg [7:0] sram_3_banks_0_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_3_banks_0_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_0_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_0_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_0_banksymbol_read_3;
  reg [7:0] sram_3_banks_1_bank_symbol0 [0:15];
  reg [7:0] sram_3_banks_1_bank_symbol1 [0:15];
  reg [7:0] sram_3_banks_1_bank_symbol2 [0:15];
  reg [7:0] sram_3_banks_1_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_3_banks_1_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_1_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_1_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_1_banksymbol_read_3;
  reg [7:0] sram_3_banks_2_bank_symbol0 [0:15];
  reg [7:0] sram_3_banks_2_bank_symbol1 [0:15];
  reg [7:0] sram_3_banks_2_bank_symbol2 [0:15];
  reg [7:0] sram_3_banks_2_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_3_banks_2_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_2_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_2_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_2_banksymbol_read_3;
  reg [7:0] sram_3_banks_3_bank_symbol0 [0:15];
  reg [7:0] sram_3_banks_3_bank_symbol1 [0:15];
  reg [7:0] sram_3_banks_3_bank_symbol2 [0:15];
  reg [7:0] sram_3_banks_3_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_3_banks_3_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_3_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_3_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_3_banksymbol_read_3;
  reg [7:0] sram_3_banks_4_bank_symbol0 [0:15];
  reg [7:0] sram_3_banks_4_bank_symbol1 [0:15];
  reg [7:0] sram_3_banks_4_bank_symbol2 [0:15];
  reg [7:0] sram_3_banks_4_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_3_banks_4_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_4_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_4_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_4_banksymbol_read_3;
  reg [7:0] sram_3_banks_5_bank_symbol0 [0:15];
  reg [7:0] sram_3_banks_5_bank_symbol1 [0:15];
  reg [7:0] sram_3_banks_5_bank_symbol2 [0:15];
  reg [7:0] sram_3_banks_5_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_3_banks_5_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_5_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_5_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_5_banksymbol_read_3;
  reg [7:0] sram_3_banks_6_bank_symbol0 [0:15];
  reg [7:0] sram_3_banks_6_bank_symbol1 [0:15];
  reg [7:0] sram_3_banks_6_bank_symbol2 [0:15];
  reg [7:0] sram_3_banks_6_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_3_banks_6_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_6_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_6_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_6_banksymbol_read_3;
  reg [7:0] sram_3_banks_7_bank_symbol0 [0:15];
  reg [7:0] sram_3_banks_7_bank_symbol1 [0:15];
  reg [7:0] sram_3_banks_7_bank_symbol2 [0:15];
  reg [7:0] sram_3_banks_7_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_3_banks_7_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_7_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_7_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_7_banksymbol_read_3;
  reg [7:0] sram_3_banks_8_bank_symbol0 [0:15];
  reg [7:0] sram_3_banks_8_bank_symbol1 [0:15];
  reg [7:0] sram_3_banks_8_bank_symbol2 [0:15];
  reg [7:0] sram_3_banks_8_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_3_banks_8_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_8_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_8_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_8_banksymbol_read_3;
  reg [7:0] sram_3_banks_9_bank_symbol0 [0:15];
  reg [7:0] sram_3_banks_9_bank_symbol1 [0:15];
  reg [7:0] sram_3_banks_9_bank_symbol2 [0:15];
  reg [7:0] sram_3_banks_9_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_3_banks_9_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_9_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_9_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_9_banksymbol_read_3;
  reg [7:0] sram_3_banks_10_bank_symbol0 [0:15];
  reg [7:0] sram_3_banks_10_bank_symbol1 [0:15];
  reg [7:0] sram_3_banks_10_bank_symbol2 [0:15];
  reg [7:0] sram_3_banks_10_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_3_banks_10_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_10_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_10_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_10_banksymbol_read_3;
  reg [7:0] sram_3_banks_11_bank_symbol0 [0:15];
  reg [7:0] sram_3_banks_11_bank_symbol1 [0:15];
  reg [7:0] sram_3_banks_11_bank_symbol2 [0:15];
  reg [7:0] sram_3_banks_11_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_3_banks_11_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_11_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_11_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_11_banksymbol_read_3;
  reg [7:0] sram_3_banks_12_bank_symbol0 [0:15];
  reg [7:0] sram_3_banks_12_bank_symbol1 [0:15];
  reg [7:0] sram_3_banks_12_bank_symbol2 [0:15];
  reg [7:0] sram_3_banks_12_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_3_banks_12_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_12_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_12_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_12_banksymbol_read_3;
  reg [7:0] sram_3_banks_13_bank_symbol0 [0:15];
  reg [7:0] sram_3_banks_13_bank_symbol1 [0:15];
  reg [7:0] sram_3_banks_13_bank_symbol2 [0:15];
  reg [7:0] sram_3_banks_13_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_3_banks_13_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_13_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_13_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_13_banksymbol_read_3;
  reg [7:0] sram_3_banks_14_bank_symbol0 [0:15];
  reg [7:0] sram_3_banks_14_bank_symbol1 [0:15];
  reg [7:0] sram_3_banks_14_bank_symbol2 [0:15];
  reg [7:0] sram_3_banks_14_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_3_banks_14_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_14_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_14_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_14_banksymbol_read_3;
  reg [7:0] sram_3_banks_15_bank_symbol0 [0:15];
  reg [7:0] sram_3_banks_15_bank_symbol1 [0:15];
  reg [7:0] sram_3_banks_15_bank_symbol2 [0:15];
  reg [7:0] sram_3_banks_15_bank_symbol3 [0:15];
  reg [7:0] _zz_sram_3_banks_15_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_15_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_15_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_15_banksymbol_read_3;

  assign _zz_sram_0_banks_0_bank_port = sram_0_ports_cmd_payload_wdata[31 : 0];
  assign _zz_sram_0_banks_0_bank_port_1 = sram_0_ports_cmd_payload_wstrb[3 : 0];
  assign _zz_sram_0_banks_0_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[0]);
  assign _zz_sram_0_banks_1_bank_port = sram_0_ports_cmd_payload_wdata[63 : 32];
  assign _zz_sram_0_banks_1_bank_port_1 = sram_0_ports_cmd_payload_wstrb[7 : 4];
  assign _zz_sram_0_banks_1_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[1]);
  assign _zz_sram_0_banks_2_bank_port = sram_0_ports_cmd_payload_wdata[95 : 64];
  assign _zz_sram_0_banks_2_bank_port_1 = sram_0_ports_cmd_payload_wstrb[11 : 8];
  assign _zz_sram_0_banks_2_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[2]);
  assign _zz_sram_0_banks_3_bank_port = sram_0_ports_cmd_payload_wdata[127 : 96];
  assign _zz_sram_0_banks_3_bank_port_1 = sram_0_ports_cmd_payload_wstrb[15 : 12];
  assign _zz_sram_0_banks_3_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[3]);
  assign _zz_sram_0_banks_4_bank_port = sram_0_ports_cmd_payload_wdata[159 : 128];
  assign _zz_sram_0_banks_4_bank_port_1 = sram_0_ports_cmd_payload_wstrb[19 : 16];
  assign _zz_sram_0_banks_4_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[4]);
  assign _zz_sram_0_banks_5_bank_port = sram_0_ports_cmd_payload_wdata[191 : 160];
  assign _zz_sram_0_banks_5_bank_port_1 = sram_0_ports_cmd_payload_wstrb[23 : 20];
  assign _zz_sram_0_banks_5_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[5]);
  assign _zz_sram_0_banks_6_bank_port = sram_0_ports_cmd_payload_wdata[223 : 192];
  assign _zz_sram_0_banks_6_bank_port_1 = sram_0_ports_cmd_payload_wstrb[27 : 24];
  assign _zz_sram_0_banks_6_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[6]);
  assign _zz_sram_0_banks_7_bank_port = sram_0_ports_cmd_payload_wdata[255 : 224];
  assign _zz_sram_0_banks_7_bank_port_1 = sram_0_ports_cmd_payload_wstrb[31 : 28];
  assign _zz_sram_0_banks_7_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[7]);
  assign _zz_sram_0_banks_8_bank_port = sram_0_ports_cmd_payload_wdata[287 : 256];
  assign _zz_sram_0_banks_8_bank_port_1 = sram_0_ports_cmd_payload_wstrb[35 : 32];
  assign _zz_sram_0_banks_8_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[8]);
  assign _zz_sram_0_banks_9_bank_port = sram_0_ports_cmd_payload_wdata[319 : 288];
  assign _zz_sram_0_banks_9_bank_port_1 = sram_0_ports_cmd_payload_wstrb[39 : 36];
  assign _zz_sram_0_banks_9_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[9]);
  assign _zz_sram_0_banks_10_bank_port = sram_0_ports_cmd_payload_wdata[351 : 320];
  assign _zz_sram_0_banks_10_bank_port_1 = sram_0_ports_cmd_payload_wstrb[43 : 40];
  assign _zz_sram_0_banks_10_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[10]);
  assign _zz_sram_0_banks_11_bank_port = sram_0_ports_cmd_payload_wdata[383 : 352];
  assign _zz_sram_0_banks_11_bank_port_1 = sram_0_ports_cmd_payload_wstrb[47 : 44];
  assign _zz_sram_0_banks_11_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[11]);
  assign _zz_sram_0_banks_12_bank_port = sram_0_ports_cmd_payload_wdata[415 : 384];
  assign _zz_sram_0_banks_12_bank_port_1 = sram_0_ports_cmd_payload_wstrb[51 : 48];
  assign _zz_sram_0_banks_12_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[12]);
  assign _zz_sram_0_banks_13_bank_port = sram_0_ports_cmd_payload_wdata[447 : 416];
  assign _zz_sram_0_banks_13_bank_port_1 = sram_0_ports_cmd_payload_wstrb[55 : 52];
  assign _zz_sram_0_banks_13_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[13]);
  assign _zz_sram_0_banks_14_bank_port = sram_0_ports_cmd_payload_wdata[479 : 448];
  assign _zz_sram_0_banks_14_bank_port_1 = sram_0_ports_cmd_payload_wstrb[59 : 56];
  assign _zz_sram_0_banks_14_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[14]);
  assign _zz_sram_0_banks_15_bank_port = sram_0_ports_cmd_payload_wdata[511 : 480];
  assign _zz_sram_0_banks_15_bank_port_1 = sram_0_ports_cmd_payload_wstrb[63 : 60];
  assign _zz_sram_0_banks_15_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[15]);
  assign _zz_sram_1_banks_0_bank_port = sram_1_ports_cmd_payload_wdata[31 : 0];
  assign _zz_sram_1_banks_0_bank_port_1 = sram_1_ports_cmd_payload_wstrb[3 : 0];
  assign _zz_sram_1_banks_0_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[0]);
  assign _zz_sram_1_banks_1_bank_port = sram_1_ports_cmd_payload_wdata[63 : 32];
  assign _zz_sram_1_banks_1_bank_port_1 = sram_1_ports_cmd_payload_wstrb[7 : 4];
  assign _zz_sram_1_banks_1_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[1]);
  assign _zz_sram_1_banks_2_bank_port = sram_1_ports_cmd_payload_wdata[95 : 64];
  assign _zz_sram_1_banks_2_bank_port_1 = sram_1_ports_cmd_payload_wstrb[11 : 8];
  assign _zz_sram_1_banks_2_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[2]);
  assign _zz_sram_1_banks_3_bank_port = sram_1_ports_cmd_payload_wdata[127 : 96];
  assign _zz_sram_1_banks_3_bank_port_1 = sram_1_ports_cmd_payload_wstrb[15 : 12];
  assign _zz_sram_1_banks_3_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[3]);
  assign _zz_sram_1_banks_4_bank_port = sram_1_ports_cmd_payload_wdata[159 : 128];
  assign _zz_sram_1_banks_4_bank_port_1 = sram_1_ports_cmd_payload_wstrb[19 : 16];
  assign _zz_sram_1_banks_4_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[4]);
  assign _zz_sram_1_banks_5_bank_port = sram_1_ports_cmd_payload_wdata[191 : 160];
  assign _zz_sram_1_banks_5_bank_port_1 = sram_1_ports_cmd_payload_wstrb[23 : 20];
  assign _zz_sram_1_banks_5_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[5]);
  assign _zz_sram_1_banks_6_bank_port = sram_1_ports_cmd_payload_wdata[223 : 192];
  assign _zz_sram_1_banks_6_bank_port_1 = sram_1_ports_cmd_payload_wstrb[27 : 24];
  assign _zz_sram_1_banks_6_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[6]);
  assign _zz_sram_1_banks_7_bank_port = sram_1_ports_cmd_payload_wdata[255 : 224];
  assign _zz_sram_1_banks_7_bank_port_1 = sram_1_ports_cmd_payload_wstrb[31 : 28];
  assign _zz_sram_1_banks_7_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[7]);
  assign _zz_sram_1_banks_8_bank_port = sram_1_ports_cmd_payload_wdata[287 : 256];
  assign _zz_sram_1_banks_8_bank_port_1 = sram_1_ports_cmd_payload_wstrb[35 : 32];
  assign _zz_sram_1_banks_8_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[8]);
  assign _zz_sram_1_banks_9_bank_port = sram_1_ports_cmd_payload_wdata[319 : 288];
  assign _zz_sram_1_banks_9_bank_port_1 = sram_1_ports_cmd_payload_wstrb[39 : 36];
  assign _zz_sram_1_banks_9_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[9]);
  assign _zz_sram_1_banks_10_bank_port = sram_1_ports_cmd_payload_wdata[351 : 320];
  assign _zz_sram_1_banks_10_bank_port_1 = sram_1_ports_cmd_payload_wstrb[43 : 40];
  assign _zz_sram_1_banks_10_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[10]);
  assign _zz_sram_1_banks_11_bank_port = sram_1_ports_cmd_payload_wdata[383 : 352];
  assign _zz_sram_1_banks_11_bank_port_1 = sram_1_ports_cmd_payload_wstrb[47 : 44];
  assign _zz_sram_1_banks_11_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[11]);
  assign _zz_sram_1_banks_12_bank_port = sram_1_ports_cmd_payload_wdata[415 : 384];
  assign _zz_sram_1_banks_12_bank_port_1 = sram_1_ports_cmd_payload_wstrb[51 : 48];
  assign _zz_sram_1_banks_12_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[12]);
  assign _zz_sram_1_banks_13_bank_port = sram_1_ports_cmd_payload_wdata[447 : 416];
  assign _zz_sram_1_banks_13_bank_port_1 = sram_1_ports_cmd_payload_wstrb[55 : 52];
  assign _zz_sram_1_banks_13_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[13]);
  assign _zz_sram_1_banks_14_bank_port = sram_1_ports_cmd_payload_wdata[479 : 448];
  assign _zz_sram_1_banks_14_bank_port_1 = sram_1_ports_cmd_payload_wstrb[59 : 56];
  assign _zz_sram_1_banks_14_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[14]);
  assign _zz_sram_1_banks_15_bank_port = sram_1_ports_cmd_payload_wdata[511 : 480];
  assign _zz_sram_1_banks_15_bank_port_1 = sram_1_ports_cmd_payload_wstrb[63 : 60];
  assign _zz_sram_1_banks_15_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[15]);
  assign _zz_sram_2_banks_0_bank_port = sram_2_ports_cmd_payload_wdata[31 : 0];
  assign _zz_sram_2_banks_0_bank_port_1 = sram_2_ports_cmd_payload_wstrb[3 : 0];
  assign _zz_sram_2_banks_0_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[0]);
  assign _zz_sram_2_banks_1_bank_port = sram_2_ports_cmd_payload_wdata[63 : 32];
  assign _zz_sram_2_banks_1_bank_port_1 = sram_2_ports_cmd_payload_wstrb[7 : 4];
  assign _zz_sram_2_banks_1_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[1]);
  assign _zz_sram_2_banks_2_bank_port = sram_2_ports_cmd_payload_wdata[95 : 64];
  assign _zz_sram_2_banks_2_bank_port_1 = sram_2_ports_cmd_payload_wstrb[11 : 8];
  assign _zz_sram_2_banks_2_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[2]);
  assign _zz_sram_2_banks_3_bank_port = sram_2_ports_cmd_payload_wdata[127 : 96];
  assign _zz_sram_2_banks_3_bank_port_1 = sram_2_ports_cmd_payload_wstrb[15 : 12];
  assign _zz_sram_2_banks_3_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[3]);
  assign _zz_sram_2_banks_4_bank_port = sram_2_ports_cmd_payload_wdata[159 : 128];
  assign _zz_sram_2_banks_4_bank_port_1 = sram_2_ports_cmd_payload_wstrb[19 : 16];
  assign _zz_sram_2_banks_4_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[4]);
  assign _zz_sram_2_banks_5_bank_port = sram_2_ports_cmd_payload_wdata[191 : 160];
  assign _zz_sram_2_banks_5_bank_port_1 = sram_2_ports_cmd_payload_wstrb[23 : 20];
  assign _zz_sram_2_banks_5_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[5]);
  assign _zz_sram_2_banks_6_bank_port = sram_2_ports_cmd_payload_wdata[223 : 192];
  assign _zz_sram_2_banks_6_bank_port_1 = sram_2_ports_cmd_payload_wstrb[27 : 24];
  assign _zz_sram_2_banks_6_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[6]);
  assign _zz_sram_2_banks_7_bank_port = sram_2_ports_cmd_payload_wdata[255 : 224];
  assign _zz_sram_2_banks_7_bank_port_1 = sram_2_ports_cmd_payload_wstrb[31 : 28];
  assign _zz_sram_2_banks_7_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[7]);
  assign _zz_sram_2_banks_8_bank_port = sram_2_ports_cmd_payload_wdata[287 : 256];
  assign _zz_sram_2_banks_8_bank_port_1 = sram_2_ports_cmd_payload_wstrb[35 : 32];
  assign _zz_sram_2_banks_8_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[8]);
  assign _zz_sram_2_banks_9_bank_port = sram_2_ports_cmd_payload_wdata[319 : 288];
  assign _zz_sram_2_banks_9_bank_port_1 = sram_2_ports_cmd_payload_wstrb[39 : 36];
  assign _zz_sram_2_banks_9_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[9]);
  assign _zz_sram_2_banks_10_bank_port = sram_2_ports_cmd_payload_wdata[351 : 320];
  assign _zz_sram_2_banks_10_bank_port_1 = sram_2_ports_cmd_payload_wstrb[43 : 40];
  assign _zz_sram_2_banks_10_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[10]);
  assign _zz_sram_2_banks_11_bank_port = sram_2_ports_cmd_payload_wdata[383 : 352];
  assign _zz_sram_2_banks_11_bank_port_1 = sram_2_ports_cmd_payload_wstrb[47 : 44];
  assign _zz_sram_2_banks_11_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[11]);
  assign _zz_sram_2_banks_12_bank_port = sram_2_ports_cmd_payload_wdata[415 : 384];
  assign _zz_sram_2_banks_12_bank_port_1 = sram_2_ports_cmd_payload_wstrb[51 : 48];
  assign _zz_sram_2_banks_12_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[12]);
  assign _zz_sram_2_banks_13_bank_port = sram_2_ports_cmd_payload_wdata[447 : 416];
  assign _zz_sram_2_banks_13_bank_port_1 = sram_2_ports_cmd_payload_wstrb[55 : 52];
  assign _zz_sram_2_banks_13_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[13]);
  assign _zz_sram_2_banks_14_bank_port = sram_2_ports_cmd_payload_wdata[479 : 448];
  assign _zz_sram_2_banks_14_bank_port_1 = sram_2_ports_cmd_payload_wstrb[59 : 56];
  assign _zz_sram_2_banks_14_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[14]);
  assign _zz_sram_2_banks_15_bank_port = sram_2_ports_cmd_payload_wdata[511 : 480];
  assign _zz_sram_2_banks_15_bank_port_1 = sram_2_ports_cmd_payload_wstrb[63 : 60];
  assign _zz_sram_2_banks_15_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[15]);
  assign _zz_sram_3_banks_0_bank_port = sram_3_ports_cmd_payload_wdata[31 : 0];
  assign _zz_sram_3_banks_0_bank_port_1 = sram_3_ports_cmd_payload_wstrb[3 : 0];
  assign _zz_sram_3_banks_0_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[0]);
  assign _zz_sram_3_banks_1_bank_port = sram_3_ports_cmd_payload_wdata[63 : 32];
  assign _zz_sram_3_banks_1_bank_port_1 = sram_3_ports_cmd_payload_wstrb[7 : 4];
  assign _zz_sram_3_banks_1_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[1]);
  assign _zz_sram_3_banks_2_bank_port = sram_3_ports_cmd_payload_wdata[95 : 64];
  assign _zz_sram_3_banks_2_bank_port_1 = sram_3_ports_cmd_payload_wstrb[11 : 8];
  assign _zz_sram_3_banks_2_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[2]);
  assign _zz_sram_3_banks_3_bank_port = sram_3_ports_cmd_payload_wdata[127 : 96];
  assign _zz_sram_3_banks_3_bank_port_1 = sram_3_ports_cmd_payload_wstrb[15 : 12];
  assign _zz_sram_3_banks_3_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[3]);
  assign _zz_sram_3_banks_4_bank_port = sram_3_ports_cmd_payload_wdata[159 : 128];
  assign _zz_sram_3_banks_4_bank_port_1 = sram_3_ports_cmd_payload_wstrb[19 : 16];
  assign _zz_sram_3_banks_4_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[4]);
  assign _zz_sram_3_banks_5_bank_port = sram_3_ports_cmd_payload_wdata[191 : 160];
  assign _zz_sram_3_banks_5_bank_port_1 = sram_3_ports_cmd_payload_wstrb[23 : 20];
  assign _zz_sram_3_banks_5_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[5]);
  assign _zz_sram_3_banks_6_bank_port = sram_3_ports_cmd_payload_wdata[223 : 192];
  assign _zz_sram_3_banks_6_bank_port_1 = sram_3_ports_cmd_payload_wstrb[27 : 24];
  assign _zz_sram_3_banks_6_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[6]);
  assign _zz_sram_3_banks_7_bank_port = sram_3_ports_cmd_payload_wdata[255 : 224];
  assign _zz_sram_3_banks_7_bank_port_1 = sram_3_ports_cmd_payload_wstrb[31 : 28];
  assign _zz_sram_3_banks_7_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[7]);
  assign _zz_sram_3_banks_8_bank_port = sram_3_ports_cmd_payload_wdata[287 : 256];
  assign _zz_sram_3_banks_8_bank_port_1 = sram_3_ports_cmd_payload_wstrb[35 : 32];
  assign _zz_sram_3_banks_8_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[8]);
  assign _zz_sram_3_banks_9_bank_port = sram_3_ports_cmd_payload_wdata[319 : 288];
  assign _zz_sram_3_banks_9_bank_port_1 = sram_3_ports_cmd_payload_wstrb[39 : 36];
  assign _zz_sram_3_banks_9_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[9]);
  assign _zz_sram_3_banks_10_bank_port = sram_3_ports_cmd_payload_wdata[351 : 320];
  assign _zz_sram_3_banks_10_bank_port_1 = sram_3_ports_cmd_payload_wstrb[43 : 40];
  assign _zz_sram_3_banks_10_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[10]);
  assign _zz_sram_3_banks_11_bank_port = sram_3_ports_cmd_payload_wdata[383 : 352];
  assign _zz_sram_3_banks_11_bank_port_1 = sram_3_ports_cmd_payload_wstrb[47 : 44];
  assign _zz_sram_3_banks_11_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[11]);
  assign _zz_sram_3_banks_12_bank_port = sram_3_ports_cmd_payload_wdata[415 : 384];
  assign _zz_sram_3_banks_12_bank_port_1 = sram_3_ports_cmd_payload_wstrb[51 : 48];
  assign _zz_sram_3_banks_12_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[12]);
  assign _zz_sram_3_banks_13_bank_port = sram_3_ports_cmd_payload_wdata[447 : 416];
  assign _zz_sram_3_banks_13_bank_port_1 = sram_3_ports_cmd_payload_wstrb[55 : 52];
  assign _zz_sram_3_banks_13_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[13]);
  assign _zz_sram_3_banks_14_bank_port = sram_3_ports_cmd_payload_wdata[479 : 448];
  assign _zz_sram_3_banks_14_bank_port_1 = sram_3_ports_cmd_payload_wstrb[59 : 56];
  assign _zz_sram_3_banks_14_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[14]);
  assign _zz_sram_3_banks_15_bank_port = sram_3_ports_cmd_payload_wdata[511 : 480];
  assign _zz_sram_3_banks_15_bank_port_1 = sram_3_ports_cmd_payload_wstrb[63 : 60];
  assign _zz_sram_3_banks_15_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[15]);
  always @(*) begin
    _zz_sram_0_banks_0_bank_port1 = {_zz_sram_0_banks_0_banksymbol_read_3, _zz_sram_0_banks_0_banksymbol_read_2, _zz_sram_0_banks_0_banksymbol_read_1, _zz_sram_0_banks_0_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_0_banks_0_bank_port_1[0] && _zz_sram_0_banks_0_bank_port_2) begin
      sram_0_banks_0_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_0_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_0_bank_port_1[1] && _zz_sram_0_banks_0_bank_port_2) begin
      sram_0_banks_0_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_0_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_0_bank_port_1[2] && _zz_sram_0_banks_0_bank_port_2) begin
      sram_0_banks_0_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_0_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_0_bank_port_1[3] && _zz_sram_0_banks_0_bank_port_2) begin
      sram_0_banks_0_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_0_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_0_banksymbol_read <= sram_0_banks_0_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_0_banksymbol_read_1 <= sram_0_banks_0_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_0_banksymbol_read_2 <= sram_0_banks_0_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_0_banksymbol_read_3 <= sram_0_banks_0_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_0_banks_1_bank_port1 = {_zz_sram_0_banks_1_banksymbol_read_3, _zz_sram_0_banks_1_banksymbol_read_2, _zz_sram_0_banks_1_banksymbol_read_1, _zz_sram_0_banks_1_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_0_banks_1_bank_port_1[0] && _zz_sram_0_banks_1_bank_port_2) begin
      sram_0_banks_1_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_1_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_1_bank_port_1[1] && _zz_sram_0_banks_1_bank_port_2) begin
      sram_0_banks_1_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_1_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_1_bank_port_1[2] && _zz_sram_0_banks_1_bank_port_2) begin
      sram_0_banks_1_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_1_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_1_bank_port_1[3] && _zz_sram_0_banks_1_bank_port_2) begin
      sram_0_banks_1_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_1_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_1_banksymbol_read <= sram_0_banks_1_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_1_banksymbol_read_1 <= sram_0_banks_1_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_1_banksymbol_read_2 <= sram_0_banks_1_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_1_banksymbol_read_3 <= sram_0_banks_1_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_0_banks_2_bank_port1 = {_zz_sram_0_banks_2_banksymbol_read_3, _zz_sram_0_banks_2_banksymbol_read_2, _zz_sram_0_banks_2_banksymbol_read_1, _zz_sram_0_banks_2_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_0_banks_2_bank_port_1[0] && _zz_sram_0_banks_2_bank_port_2) begin
      sram_0_banks_2_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_2_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_2_bank_port_1[1] && _zz_sram_0_banks_2_bank_port_2) begin
      sram_0_banks_2_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_2_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_2_bank_port_1[2] && _zz_sram_0_banks_2_bank_port_2) begin
      sram_0_banks_2_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_2_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_2_bank_port_1[3] && _zz_sram_0_banks_2_bank_port_2) begin
      sram_0_banks_2_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_2_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_2_banksymbol_read <= sram_0_banks_2_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_2_banksymbol_read_1 <= sram_0_banks_2_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_2_banksymbol_read_2 <= sram_0_banks_2_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_2_banksymbol_read_3 <= sram_0_banks_2_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_0_banks_3_bank_port1 = {_zz_sram_0_banks_3_banksymbol_read_3, _zz_sram_0_banks_3_banksymbol_read_2, _zz_sram_0_banks_3_banksymbol_read_1, _zz_sram_0_banks_3_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_0_banks_3_bank_port_1[0] && _zz_sram_0_banks_3_bank_port_2) begin
      sram_0_banks_3_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_3_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_3_bank_port_1[1] && _zz_sram_0_banks_3_bank_port_2) begin
      sram_0_banks_3_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_3_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_3_bank_port_1[2] && _zz_sram_0_banks_3_bank_port_2) begin
      sram_0_banks_3_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_3_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_3_bank_port_1[3] && _zz_sram_0_banks_3_bank_port_2) begin
      sram_0_banks_3_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_3_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_3_banksymbol_read <= sram_0_banks_3_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_3_banksymbol_read_1 <= sram_0_banks_3_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_3_banksymbol_read_2 <= sram_0_banks_3_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_3_banksymbol_read_3 <= sram_0_banks_3_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_0_banks_4_bank_port1 = {_zz_sram_0_banks_4_banksymbol_read_3, _zz_sram_0_banks_4_banksymbol_read_2, _zz_sram_0_banks_4_banksymbol_read_1, _zz_sram_0_banks_4_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_0_banks_4_bank_port_1[0] && _zz_sram_0_banks_4_bank_port_2) begin
      sram_0_banks_4_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_4_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_4_bank_port_1[1] && _zz_sram_0_banks_4_bank_port_2) begin
      sram_0_banks_4_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_4_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_4_bank_port_1[2] && _zz_sram_0_banks_4_bank_port_2) begin
      sram_0_banks_4_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_4_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_4_bank_port_1[3] && _zz_sram_0_banks_4_bank_port_2) begin
      sram_0_banks_4_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_4_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_4_banksymbol_read <= sram_0_banks_4_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_4_banksymbol_read_1 <= sram_0_banks_4_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_4_banksymbol_read_2 <= sram_0_banks_4_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_4_banksymbol_read_3 <= sram_0_banks_4_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_0_banks_5_bank_port1 = {_zz_sram_0_banks_5_banksymbol_read_3, _zz_sram_0_banks_5_banksymbol_read_2, _zz_sram_0_banks_5_banksymbol_read_1, _zz_sram_0_banks_5_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_0_banks_5_bank_port_1[0] && _zz_sram_0_banks_5_bank_port_2) begin
      sram_0_banks_5_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_5_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_5_bank_port_1[1] && _zz_sram_0_banks_5_bank_port_2) begin
      sram_0_banks_5_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_5_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_5_bank_port_1[2] && _zz_sram_0_banks_5_bank_port_2) begin
      sram_0_banks_5_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_5_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_5_bank_port_1[3] && _zz_sram_0_banks_5_bank_port_2) begin
      sram_0_banks_5_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_5_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_5_banksymbol_read <= sram_0_banks_5_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_5_banksymbol_read_1 <= sram_0_banks_5_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_5_banksymbol_read_2 <= sram_0_banks_5_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_5_banksymbol_read_3 <= sram_0_banks_5_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_0_banks_6_bank_port1 = {_zz_sram_0_banks_6_banksymbol_read_3, _zz_sram_0_banks_6_banksymbol_read_2, _zz_sram_0_banks_6_banksymbol_read_1, _zz_sram_0_banks_6_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_0_banks_6_bank_port_1[0] && _zz_sram_0_banks_6_bank_port_2) begin
      sram_0_banks_6_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_6_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_6_bank_port_1[1] && _zz_sram_0_banks_6_bank_port_2) begin
      sram_0_banks_6_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_6_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_6_bank_port_1[2] && _zz_sram_0_banks_6_bank_port_2) begin
      sram_0_banks_6_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_6_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_6_bank_port_1[3] && _zz_sram_0_banks_6_bank_port_2) begin
      sram_0_banks_6_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_6_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_6_banksymbol_read <= sram_0_banks_6_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_6_banksymbol_read_1 <= sram_0_banks_6_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_6_banksymbol_read_2 <= sram_0_banks_6_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_6_banksymbol_read_3 <= sram_0_banks_6_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_0_banks_7_bank_port1 = {_zz_sram_0_banks_7_banksymbol_read_3, _zz_sram_0_banks_7_banksymbol_read_2, _zz_sram_0_banks_7_banksymbol_read_1, _zz_sram_0_banks_7_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_0_banks_7_bank_port_1[0] && _zz_sram_0_banks_7_bank_port_2) begin
      sram_0_banks_7_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_7_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_7_bank_port_1[1] && _zz_sram_0_banks_7_bank_port_2) begin
      sram_0_banks_7_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_7_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_7_bank_port_1[2] && _zz_sram_0_banks_7_bank_port_2) begin
      sram_0_banks_7_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_7_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_7_bank_port_1[3] && _zz_sram_0_banks_7_bank_port_2) begin
      sram_0_banks_7_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_7_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_7_banksymbol_read <= sram_0_banks_7_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_7_banksymbol_read_1 <= sram_0_banks_7_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_7_banksymbol_read_2 <= sram_0_banks_7_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_7_banksymbol_read_3 <= sram_0_banks_7_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_0_banks_8_bank_port1 = {_zz_sram_0_banks_8_banksymbol_read_3, _zz_sram_0_banks_8_banksymbol_read_2, _zz_sram_0_banks_8_banksymbol_read_1, _zz_sram_0_banks_8_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_0_banks_8_bank_port_1[0] && _zz_sram_0_banks_8_bank_port_2) begin
      sram_0_banks_8_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_8_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_8_bank_port_1[1] && _zz_sram_0_banks_8_bank_port_2) begin
      sram_0_banks_8_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_8_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_8_bank_port_1[2] && _zz_sram_0_banks_8_bank_port_2) begin
      sram_0_banks_8_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_8_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_8_bank_port_1[3] && _zz_sram_0_banks_8_bank_port_2) begin
      sram_0_banks_8_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_8_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_8_banksymbol_read <= sram_0_banks_8_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_8_banksymbol_read_1 <= sram_0_banks_8_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_8_banksymbol_read_2 <= sram_0_banks_8_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_8_banksymbol_read_3 <= sram_0_banks_8_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_0_banks_9_bank_port1 = {_zz_sram_0_banks_9_banksymbol_read_3, _zz_sram_0_banks_9_banksymbol_read_2, _zz_sram_0_banks_9_banksymbol_read_1, _zz_sram_0_banks_9_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_0_banks_9_bank_port_1[0] && _zz_sram_0_banks_9_bank_port_2) begin
      sram_0_banks_9_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_9_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_9_bank_port_1[1] && _zz_sram_0_banks_9_bank_port_2) begin
      sram_0_banks_9_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_9_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_9_bank_port_1[2] && _zz_sram_0_banks_9_bank_port_2) begin
      sram_0_banks_9_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_9_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_9_bank_port_1[3] && _zz_sram_0_banks_9_bank_port_2) begin
      sram_0_banks_9_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_9_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_9_banksymbol_read <= sram_0_banks_9_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_9_banksymbol_read_1 <= sram_0_banks_9_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_9_banksymbol_read_2 <= sram_0_banks_9_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_9_banksymbol_read_3 <= sram_0_banks_9_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_0_banks_10_bank_port1 = {_zz_sram_0_banks_10_banksymbol_read_3, _zz_sram_0_banks_10_banksymbol_read_2, _zz_sram_0_banks_10_banksymbol_read_1, _zz_sram_0_banks_10_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_0_banks_10_bank_port_1[0] && _zz_sram_0_banks_10_bank_port_2) begin
      sram_0_banks_10_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_10_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_10_bank_port_1[1] && _zz_sram_0_banks_10_bank_port_2) begin
      sram_0_banks_10_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_10_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_10_bank_port_1[2] && _zz_sram_0_banks_10_bank_port_2) begin
      sram_0_banks_10_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_10_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_10_bank_port_1[3] && _zz_sram_0_banks_10_bank_port_2) begin
      sram_0_banks_10_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_10_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_10_banksymbol_read <= sram_0_banks_10_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_10_banksymbol_read_1 <= sram_0_banks_10_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_10_banksymbol_read_2 <= sram_0_banks_10_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_10_banksymbol_read_3 <= sram_0_banks_10_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_0_banks_11_bank_port1 = {_zz_sram_0_banks_11_banksymbol_read_3, _zz_sram_0_banks_11_banksymbol_read_2, _zz_sram_0_banks_11_banksymbol_read_1, _zz_sram_0_banks_11_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_0_banks_11_bank_port_1[0] && _zz_sram_0_banks_11_bank_port_2) begin
      sram_0_banks_11_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_11_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_11_bank_port_1[1] && _zz_sram_0_banks_11_bank_port_2) begin
      sram_0_banks_11_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_11_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_11_bank_port_1[2] && _zz_sram_0_banks_11_bank_port_2) begin
      sram_0_banks_11_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_11_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_11_bank_port_1[3] && _zz_sram_0_banks_11_bank_port_2) begin
      sram_0_banks_11_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_11_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_11_banksymbol_read <= sram_0_banks_11_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_11_banksymbol_read_1 <= sram_0_banks_11_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_11_banksymbol_read_2 <= sram_0_banks_11_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_11_banksymbol_read_3 <= sram_0_banks_11_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_0_banks_12_bank_port1 = {_zz_sram_0_banks_12_banksymbol_read_3, _zz_sram_0_banks_12_banksymbol_read_2, _zz_sram_0_banks_12_banksymbol_read_1, _zz_sram_0_banks_12_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_0_banks_12_bank_port_1[0] && _zz_sram_0_banks_12_bank_port_2) begin
      sram_0_banks_12_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_12_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_12_bank_port_1[1] && _zz_sram_0_banks_12_bank_port_2) begin
      sram_0_banks_12_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_12_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_12_bank_port_1[2] && _zz_sram_0_banks_12_bank_port_2) begin
      sram_0_banks_12_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_12_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_12_bank_port_1[3] && _zz_sram_0_banks_12_bank_port_2) begin
      sram_0_banks_12_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_12_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_12_banksymbol_read <= sram_0_banks_12_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_12_banksymbol_read_1 <= sram_0_banks_12_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_12_banksymbol_read_2 <= sram_0_banks_12_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_12_banksymbol_read_3 <= sram_0_banks_12_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_0_banks_13_bank_port1 = {_zz_sram_0_banks_13_banksymbol_read_3, _zz_sram_0_banks_13_banksymbol_read_2, _zz_sram_0_banks_13_banksymbol_read_1, _zz_sram_0_banks_13_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_0_banks_13_bank_port_1[0] && _zz_sram_0_banks_13_bank_port_2) begin
      sram_0_banks_13_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_13_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_13_bank_port_1[1] && _zz_sram_0_banks_13_bank_port_2) begin
      sram_0_banks_13_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_13_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_13_bank_port_1[2] && _zz_sram_0_banks_13_bank_port_2) begin
      sram_0_banks_13_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_13_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_13_bank_port_1[3] && _zz_sram_0_banks_13_bank_port_2) begin
      sram_0_banks_13_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_13_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_13_banksymbol_read <= sram_0_banks_13_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_13_banksymbol_read_1 <= sram_0_banks_13_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_13_banksymbol_read_2 <= sram_0_banks_13_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_13_banksymbol_read_3 <= sram_0_banks_13_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_0_banks_14_bank_port1 = {_zz_sram_0_banks_14_banksymbol_read_3, _zz_sram_0_banks_14_banksymbol_read_2, _zz_sram_0_banks_14_banksymbol_read_1, _zz_sram_0_banks_14_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_0_banks_14_bank_port_1[0] && _zz_sram_0_banks_14_bank_port_2) begin
      sram_0_banks_14_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_14_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_14_bank_port_1[1] && _zz_sram_0_banks_14_bank_port_2) begin
      sram_0_banks_14_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_14_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_14_bank_port_1[2] && _zz_sram_0_banks_14_bank_port_2) begin
      sram_0_banks_14_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_14_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_14_bank_port_1[3] && _zz_sram_0_banks_14_bank_port_2) begin
      sram_0_banks_14_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_14_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_14_banksymbol_read <= sram_0_banks_14_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_14_banksymbol_read_1 <= sram_0_banks_14_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_14_banksymbol_read_2 <= sram_0_banks_14_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_14_banksymbol_read_3 <= sram_0_banks_14_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_0_banks_15_bank_port1 = {_zz_sram_0_banks_15_banksymbol_read_3, _zz_sram_0_banks_15_banksymbol_read_2, _zz_sram_0_banks_15_banksymbol_read_1, _zz_sram_0_banks_15_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_0_banks_15_bank_port_1[0] && _zz_sram_0_banks_15_bank_port_2) begin
      sram_0_banks_15_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_15_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_15_bank_port_1[1] && _zz_sram_0_banks_15_bank_port_2) begin
      sram_0_banks_15_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_15_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_15_bank_port_1[2] && _zz_sram_0_banks_15_bank_port_2) begin
      sram_0_banks_15_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_15_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_15_bank_port_1[3] && _zz_sram_0_banks_15_bank_port_2) begin
      sram_0_banks_15_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_15_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_15_banksymbol_read <= sram_0_banks_15_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_15_banksymbol_read_1 <= sram_0_banks_15_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_15_banksymbol_read_2 <= sram_0_banks_15_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_15_banksymbol_read_3 <= sram_0_banks_15_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_0_bank_port1 = {_zz_sram_1_banks_0_banksymbol_read_3, _zz_sram_1_banks_0_banksymbol_read_2, _zz_sram_1_banks_0_banksymbol_read_1, _zz_sram_1_banks_0_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_1_banks_0_bank_port_1[0] && _zz_sram_1_banks_0_bank_port_2) begin
      sram_1_banks_0_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_0_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_0_bank_port_1[1] && _zz_sram_1_banks_0_bank_port_2) begin
      sram_1_banks_0_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_0_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_0_bank_port_1[2] && _zz_sram_1_banks_0_bank_port_2) begin
      sram_1_banks_0_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_0_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_0_bank_port_1[3] && _zz_sram_1_banks_0_bank_port_2) begin
      sram_1_banks_0_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_0_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_0_banksymbol_read <= sram_1_banks_0_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_0_banksymbol_read_1 <= sram_1_banks_0_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_0_banksymbol_read_2 <= sram_1_banks_0_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_0_banksymbol_read_3 <= sram_1_banks_0_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_1_bank_port1 = {_zz_sram_1_banks_1_banksymbol_read_3, _zz_sram_1_banks_1_banksymbol_read_2, _zz_sram_1_banks_1_banksymbol_read_1, _zz_sram_1_banks_1_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_1_banks_1_bank_port_1[0] && _zz_sram_1_banks_1_bank_port_2) begin
      sram_1_banks_1_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_1_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_1_bank_port_1[1] && _zz_sram_1_banks_1_bank_port_2) begin
      sram_1_banks_1_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_1_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_1_bank_port_1[2] && _zz_sram_1_banks_1_bank_port_2) begin
      sram_1_banks_1_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_1_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_1_bank_port_1[3] && _zz_sram_1_banks_1_bank_port_2) begin
      sram_1_banks_1_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_1_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_1_banksymbol_read <= sram_1_banks_1_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_1_banksymbol_read_1 <= sram_1_banks_1_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_1_banksymbol_read_2 <= sram_1_banks_1_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_1_banksymbol_read_3 <= sram_1_banks_1_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_2_bank_port1 = {_zz_sram_1_banks_2_banksymbol_read_3, _zz_sram_1_banks_2_banksymbol_read_2, _zz_sram_1_banks_2_banksymbol_read_1, _zz_sram_1_banks_2_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_1_banks_2_bank_port_1[0] && _zz_sram_1_banks_2_bank_port_2) begin
      sram_1_banks_2_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_2_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_2_bank_port_1[1] && _zz_sram_1_banks_2_bank_port_2) begin
      sram_1_banks_2_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_2_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_2_bank_port_1[2] && _zz_sram_1_banks_2_bank_port_2) begin
      sram_1_banks_2_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_2_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_2_bank_port_1[3] && _zz_sram_1_banks_2_bank_port_2) begin
      sram_1_banks_2_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_2_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_2_banksymbol_read <= sram_1_banks_2_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_2_banksymbol_read_1 <= sram_1_banks_2_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_2_banksymbol_read_2 <= sram_1_banks_2_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_2_banksymbol_read_3 <= sram_1_banks_2_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_3_bank_port1 = {_zz_sram_1_banks_3_banksymbol_read_3, _zz_sram_1_banks_3_banksymbol_read_2, _zz_sram_1_banks_3_banksymbol_read_1, _zz_sram_1_banks_3_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_1_banks_3_bank_port_1[0] && _zz_sram_1_banks_3_bank_port_2) begin
      sram_1_banks_3_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_3_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_3_bank_port_1[1] && _zz_sram_1_banks_3_bank_port_2) begin
      sram_1_banks_3_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_3_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_3_bank_port_1[2] && _zz_sram_1_banks_3_bank_port_2) begin
      sram_1_banks_3_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_3_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_3_bank_port_1[3] && _zz_sram_1_banks_3_bank_port_2) begin
      sram_1_banks_3_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_3_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_3_banksymbol_read <= sram_1_banks_3_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_3_banksymbol_read_1 <= sram_1_banks_3_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_3_banksymbol_read_2 <= sram_1_banks_3_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_3_banksymbol_read_3 <= sram_1_banks_3_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_4_bank_port1 = {_zz_sram_1_banks_4_banksymbol_read_3, _zz_sram_1_banks_4_banksymbol_read_2, _zz_sram_1_banks_4_banksymbol_read_1, _zz_sram_1_banks_4_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_1_banks_4_bank_port_1[0] && _zz_sram_1_banks_4_bank_port_2) begin
      sram_1_banks_4_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_4_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_4_bank_port_1[1] && _zz_sram_1_banks_4_bank_port_2) begin
      sram_1_banks_4_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_4_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_4_bank_port_1[2] && _zz_sram_1_banks_4_bank_port_2) begin
      sram_1_banks_4_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_4_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_4_bank_port_1[3] && _zz_sram_1_banks_4_bank_port_2) begin
      sram_1_banks_4_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_4_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_4_banksymbol_read <= sram_1_banks_4_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_4_banksymbol_read_1 <= sram_1_banks_4_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_4_banksymbol_read_2 <= sram_1_banks_4_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_4_banksymbol_read_3 <= sram_1_banks_4_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_5_bank_port1 = {_zz_sram_1_banks_5_banksymbol_read_3, _zz_sram_1_banks_5_banksymbol_read_2, _zz_sram_1_banks_5_banksymbol_read_1, _zz_sram_1_banks_5_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_1_banks_5_bank_port_1[0] && _zz_sram_1_banks_5_bank_port_2) begin
      sram_1_banks_5_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_5_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_5_bank_port_1[1] && _zz_sram_1_banks_5_bank_port_2) begin
      sram_1_banks_5_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_5_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_5_bank_port_1[2] && _zz_sram_1_banks_5_bank_port_2) begin
      sram_1_banks_5_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_5_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_5_bank_port_1[3] && _zz_sram_1_banks_5_bank_port_2) begin
      sram_1_banks_5_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_5_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_5_banksymbol_read <= sram_1_banks_5_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_5_banksymbol_read_1 <= sram_1_banks_5_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_5_banksymbol_read_2 <= sram_1_banks_5_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_5_banksymbol_read_3 <= sram_1_banks_5_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_6_bank_port1 = {_zz_sram_1_banks_6_banksymbol_read_3, _zz_sram_1_banks_6_banksymbol_read_2, _zz_sram_1_banks_6_banksymbol_read_1, _zz_sram_1_banks_6_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_1_banks_6_bank_port_1[0] && _zz_sram_1_banks_6_bank_port_2) begin
      sram_1_banks_6_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_6_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_6_bank_port_1[1] && _zz_sram_1_banks_6_bank_port_2) begin
      sram_1_banks_6_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_6_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_6_bank_port_1[2] && _zz_sram_1_banks_6_bank_port_2) begin
      sram_1_banks_6_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_6_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_6_bank_port_1[3] && _zz_sram_1_banks_6_bank_port_2) begin
      sram_1_banks_6_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_6_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_6_banksymbol_read <= sram_1_banks_6_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_6_banksymbol_read_1 <= sram_1_banks_6_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_6_banksymbol_read_2 <= sram_1_banks_6_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_6_banksymbol_read_3 <= sram_1_banks_6_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_7_bank_port1 = {_zz_sram_1_banks_7_banksymbol_read_3, _zz_sram_1_banks_7_banksymbol_read_2, _zz_sram_1_banks_7_banksymbol_read_1, _zz_sram_1_banks_7_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_1_banks_7_bank_port_1[0] && _zz_sram_1_banks_7_bank_port_2) begin
      sram_1_banks_7_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_7_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_7_bank_port_1[1] && _zz_sram_1_banks_7_bank_port_2) begin
      sram_1_banks_7_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_7_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_7_bank_port_1[2] && _zz_sram_1_banks_7_bank_port_2) begin
      sram_1_banks_7_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_7_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_7_bank_port_1[3] && _zz_sram_1_banks_7_bank_port_2) begin
      sram_1_banks_7_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_7_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_7_banksymbol_read <= sram_1_banks_7_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_7_banksymbol_read_1 <= sram_1_banks_7_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_7_banksymbol_read_2 <= sram_1_banks_7_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_7_banksymbol_read_3 <= sram_1_banks_7_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_8_bank_port1 = {_zz_sram_1_banks_8_banksymbol_read_3, _zz_sram_1_banks_8_banksymbol_read_2, _zz_sram_1_banks_8_banksymbol_read_1, _zz_sram_1_banks_8_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_1_banks_8_bank_port_1[0] && _zz_sram_1_banks_8_bank_port_2) begin
      sram_1_banks_8_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_8_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_8_bank_port_1[1] && _zz_sram_1_banks_8_bank_port_2) begin
      sram_1_banks_8_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_8_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_8_bank_port_1[2] && _zz_sram_1_banks_8_bank_port_2) begin
      sram_1_banks_8_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_8_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_8_bank_port_1[3] && _zz_sram_1_banks_8_bank_port_2) begin
      sram_1_banks_8_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_8_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_8_banksymbol_read <= sram_1_banks_8_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_8_banksymbol_read_1 <= sram_1_banks_8_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_8_banksymbol_read_2 <= sram_1_banks_8_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_8_banksymbol_read_3 <= sram_1_banks_8_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_9_bank_port1 = {_zz_sram_1_banks_9_banksymbol_read_3, _zz_sram_1_banks_9_banksymbol_read_2, _zz_sram_1_banks_9_banksymbol_read_1, _zz_sram_1_banks_9_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_1_banks_9_bank_port_1[0] && _zz_sram_1_banks_9_bank_port_2) begin
      sram_1_banks_9_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_9_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_9_bank_port_1[1] && _zz_sram_1_banks_9_bank_port_2) begin
      sram_1_banks_9_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_9_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_9_bank_port_1[2] && _zz_sram_1_banks_9_bank_port_2) begin
      sram_1_banks_9_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_9_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_9_bank_port_1[3] && _zz_sram_1_banks_9_bank_port_2) begin
      sram_1_banks_9_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_9_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_9_banksymbol_read <= sram_1_banks_9_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_9_banksymbol_read_1 <= sram_1_banks_9_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_9_banksymbol_read_2 <= sram_1_banks_9_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_9_banksymbol_read_3 <= sram_1_banks_9_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_10_bank_port1 = {_zz_sram_1_banks_10_banksymbol_read_3, _zz_sram_1_banks_10_banksymbol_read_2, _zz_sram_1_banks_10_banksymbol_read_1, _zz_sram_1_banks_10_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_1_banks_10_bank_port_1[0] && _zz_sram_1_banks_10_bank_port_2) begin
      sram_1_banks_10_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_10_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_10_bank_port_1[1] && _zz_sram_1_banks_10_bank_port_2) begin
      sram_1_banks_10_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_10_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_10_bank_port_1[2] && _zz_sram_1_banks_10_bank_port_2) begin
      sram_1_banks_10_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_10_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_10_bank_port_1[3] && _zz_sram_1_banks_10_bank_port_2) begin
      sram_1_banks_10_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_10_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_10_banksymbol_read <= sram_1_banks_10_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_10_banksymbol_read_1 <= sram_1_banks_10_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_10_banksymbol_read_2 <= sram_1_banks_10_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_10_banksymbol_read_3 <= sram_1_banks_10_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_11_bank_port1 = {_zz_sram_1_banks_11_banksymbol_read_3, _zz_sram_1_banks_11_banksymbol_read_2, _zz_sram_1_banks_11_banksymbol_read_1, _zz_sram_1_banks_11_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_1_banks_11_bank_port_1[0] && _zz_sram_1_banks_11_bank_port_2) begin
      sram_1_banks_11_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_11_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_11_bank_port_1[1] && _zz_sram_1_banks_11_bank_port_2) begin
      sram_1_banks_11_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_11_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_11_bank_port_1[2] && _zz_sram_1_banks_11_bank_port_2) begin
      sram_1_banks_11_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_11_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_11_bank_port_1[3] && _zz_sram_1_banks_11_bank_port_2) begin
      sram_1_banks_11_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_11_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_11_banksymbol_read <= sram_1_banks_11_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_11_banksymbol_read_1 <= sram_1_banks_11_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_11_banksymbol_read_2 <= sram_1_banks_11_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_11_banksymbol_read_3 <= sram_1_banks_11_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_12_bank_port1 = {_zz_sram_1_banks_12_banksymbol_read_3, _zz_sram_1_banks_12_banksymbol_read_2, _zz_sram_1_banks_12_banksymbol_read_1, _zz_sram_1_banks_12_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_1_banks_12_bank_port_1[0] && _zz_sram_1_banks_12_bank_port_2) begin
      sram_1_banks_12_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_12_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_12_bank_port_1[1] && _zz_sram_1_banks_12_bank_port_2) begin
      sram_1_banks_12_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_12_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_12_bank_port_1[2] && _zz_sram_1_banks_12_bank_port_2) begin
      sram_1_banks_12_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_12_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_12_bank_port_1[3] && _zz_sram_1_banks_12_bank_port_2) begin
      sram_1_banks_12_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_12_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_12_banksymbol_read <= sram_1_banks_12_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_12_banksymbol_read_1 <= sram_1_banks_12_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_12_banksymbol_read_2 <= sram_1_banks_12_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_12_banksymbol_read_3 <= sram_1_banks_12_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_13_bank_port1 = {_zz_sram_1_banks_13_banksymbol_read_3, _zz_sram_1_banks_13_banksymbol_read_2, _zz_sram_1_banks_13_banksymbol_read_1, _zz_sram_1_banks_13_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_1_banks_13_bank_port_1[0] && _zz_sram_1_banks_13_bank_port_2) begin
      sram_1_banks_13_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_13_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_13_bank_port_1[1] && _zz_sram_1_banks_13_bank_port_2) begin
      sram_1_banks_13_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_13_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_13_bank_port_1[2] && _zz_sram_1_banks_13_bank_port_2) begin
      sram_1_banks_13_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_13_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_13_bank_port_1[3] && _zz_sram_1_banks_13_bank_port_2) begin
      sram_1_banks_13_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_13_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_13_banksymbol_read <= sram_1_banks_13_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_13_banksymbol_read_1 <= sram_1_banks_13_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_13_banksymbol_read_2 <= sram_1_banks_13_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_13_banksymbol_read_3 <= sram_1_banks_13_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_14_bank_port1 = {_zz_sram_1_banks_14_banksymbol_read_3, _zz_sram_1_banks_14_banksymbol_read_2, _zz_sram_1_banks_14_banksymbol_read_1, _zz_sram_1_banks_14_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_1_banks_14_bank_port_1[0] && _zz_sram_1_banks_14_bank_port_2) begin
      sram_1_banks_14_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_14_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_14_bank_port_1[1] && _zz_sram_1_banks_14_bank_port_2) begin
      sram_1_banks_14_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_14_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_14_bank_port_1[2] && _zz_sram_1_banks_14_bank_port_2) begin
      sram_1_banks_14_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_14_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_14_bank_port_1[3] && _zz_sram_1_banks_14_bank_port_2) begin
      sram_1_banks_14_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_14_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_14_banksymbol_read <= sram_1_banks_14_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_14_banksymbol_read_1 <= sram_1_banks_14_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_14_banksymbol_read_2 <= sram_1_banks_14_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_14_banksymbol_read_3 <= sram_1_banks_14_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_15_bank_port1 = {_zz_sram_1_banks_15_banksymbol_read_3, _zz_sram_1_banks_15_banksymbol_read_2, _zz_sram_1_banks_15_banksymbol_read_1, _zz_sram_1_banks_15_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_1_banks_15_bank_port_1[0] && _zz_sram_1_banks_15_bank_port_2) begin
      sram_1_banks_15_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_15_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_15_bank_port_1[1] && _zz_sram_1_banks_15_bank_port_2) begin
      sram_1_banks_15_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_15_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_15_bank_port_1[2] && _zz_sram_1_banks_15_bank_port_2) begin
      sram_1_banks_15_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_15_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_15_bank_port_1[3] && _zz_sram_1_banks_15_bank_port_2) begin
      sram_1_banks_15_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_15_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_15_banksymbol_read <= sram_1_banks_15_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_15_banksymbol_read_1 <= sram_1_banks_15_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_15_banksymbol_read_2 <= sram_1_banks_15_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_15_banksymbol_read_3 <= sram_1_banks_15_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_0_bank_port1 = {_zz_sram_2_banks_0_banksymbol_read_3, _zz_sram_2_banks_0_banksymbol_read_2, _zz_sram_2_banks_0_banksymbol_read_1, _zz_sram_2_banks_0_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_2_banks_0_bank_port_1[0] && _zz_sram_2_banks_0_bank_port_2) begin
      sram_2_banks_0_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_0_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_0_bank_port_1[1] && _zz_sram_2_banks_0_bank_port_2) begin
      sram_2_banks_0_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_0_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_0_bank_port_1[2] && _zz_sram_2_banks_0_bank_port_2) begin
      sram_2_banks_0_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_0_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_0_bank_port_1[3] && _zz_sram_2_banks_0_bank_port_2) begin
      sram_2_banks_0_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_0_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_0_banksymbol_read <= sram_2_banks_0_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_0_banksymbol_read_1 <= sram_2_banks_0_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_0_banksymbol_read_2 <= sram_2_banks_0_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_0_banksymbol_read_3 <= sram_2_banks_0_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_1_bank_port1 = {_zz_sram_2_banks_1_banksymbol_read_3, _zz_sram_2_banks_1_banksymbol_read_2, _zz_sram_2_banks_1_banksymbol_read_1, _zz_sram_2_banks_1_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_2_banks_1_bank_port_1[0] && _zz_sram_2_banks_1_bank_port_2) begin
      sram_2_banks_1_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_1_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_1_bank_port_1[1] && _zz_sram_2_banks_1_bank_port_2) begin
      sram_2_banks_1_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_1_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_1_bank_port_1[2] && _zz_sram_2_banks_1_bank_port_2) begin
      sram_2_banks_1_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_1_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_1_bank_port_1[3] && _zz_sram_2_banks_1_bank_port_2) begin
      sram_2_banks_1_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_1_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_1_banksymbol_read <= sram_2_banks_1_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_1_banksymbol_read_1 <= sram_2_banks_1_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_1_banksymbol_read_2 <= sram_2_banks_1_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_1_banksymbol_read_3 <= sram_2_banks_1_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_2_bank_port1 = {_zz_sram_2_banks_2_banksymbol_read_3, _zz_sram_2_banks_2_banksymbol_read_2, _zz_sram_2_banks_2_banksymbol_read_1, _zz_sram_2_banks_2_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_2_banks_2_bank_port_1[0] && _zz_sram_2_banks_2_bank_port_2) begin
      sram_2_banks_2_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_2_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_2_bank_port_1[1] && _zz_sram_2_banks_2_bank_port_2) begin
      sram_2_banks_2_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_2_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_2_bank_port_1[2] && _zz_sram_2_banks_2_bank_port_2) begin
      sram_2_banks_2_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_2_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_2_bank_port_1[3] && _zz_sram_2_banks_2_bank_port_2) begin
      sram_2_banks_2_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_2_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_2_banksymbol_read <= sram_2_banks_2_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_2_banksymbol_read_1 <= sram_2_banks_2_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_2_banksymbol_read_2 <= sram_2_banks_2_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_2_banksymbol_read_3 <= sram_2_banks_2_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_3_bank_port1 = {_zz_sram_2_banks_3_banksymbol_read_3, _zz_sram_2_banks_3_banksymbol_read_2, _zz_sram_2_banks_3_banksymbol_read_1, _zz_sram_2_banks_3_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_2_banks_3_bank_port_1[0] && _zz_sram_2_banks_3_bank_port_2) begin
      sram_2_banks_3_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_3_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_3_bank_port_1[1] && _zz_sram_2_banks_3_bank_port_2) begin
      sram_2_banks_3_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_3_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_3_bank_port_1[2] && _zz_sram_2_banks_3_bank_port_2) begin
      sram_2_banks_3_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_3_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_3_bank_port_1[3] && _zz_sram_2_banks_3_bank_port_2) begin
      sram_2_banks_3_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_3_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_3_banksymbol_read <= sram_2_banks_3_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_3_banksymbol_read_1 <= sram_2_banks_3_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_3_banksymbol_read_2 <= sram_2_banks_3_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_3_banksymbol_read_3 <= sram_2_banks_3_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_4_bank_port1 = {_zz_sram_2_banks_4_banksymbol_read_3, _zz_sram_2_banks_4_banksymbol_read_2, _zz_sram_2_banks_4_banksymbol_read_1, _zz_sram_2_banks_4_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_2_banks_4_bank_port_1[0] && _zz_sram_2_banks_4_bank_port_2) begin
      sram_2_banks_4_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_4_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_4_bank_port_1[1] && _zz_sram_2_banks_4_bank_port_2) begin
      sram_2_banks_4_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_4_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_4_bank_port_1[2] && _zz_sram_2_banks_4_bank_port_2) begin
      sram_2_banks_4_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_4_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_4_bank_port_1[3] && _zz_sram_2_banks_4_bank_port_2) begin
      sram_2_banks_4_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_4_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_4_banksymbol_read <= sram_2_banks_4_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_4_banksymbol_read_1 <= sram_2_banks_4_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_4_banksymbol_read_2 <= sram_2_banks_4_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_4_banksymbol_read_3 <= sram_2_banks_4_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_5_bank_port1 = {_zz_sram_2_banks_5_banksymbol_read_3, _zz_sram_2_banks_5_banksymbol_read_2, _zz_sram_2_banks_5_banksymbol_read_1, _zz_sram_2_banks_5_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_2_banks_5_bank_port_1[0] && _zz_sram_2_banks_5_bank_port_2) begin
      sram_2_banks_5_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_5_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_5_bank_port_1[1] && _zz_sram_2_banks_5_bank_port_2) begin
      sram_2_banks_5_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_5_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_5_bank_port_1[2] && _zz_sram_2_banks_5_bank_port_2) begin
      sram_2_banks_5_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_5_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_5_bank_port_1[3] && _zz_sram_2_banks_5_bank_port_2) begin
      sram_2_banks_5_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_5_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_5_banksymbol_read <= sram_2_banks_5_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_5_banksymbol_read_1 <= sram_2_banks_5_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_5_banksymbol_read_2 <= sram_2_banks_5_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_5_banksymbol_read_3 <= sram_2_banks_5_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_6_bank_port1 = {_zz_sram_2_banks_6_banksymbol_read_3, _zz_sram_2_banks_6_banksymbol_read_2, _zz_sram_2_banks_6_banksymbol_read_1, _zz_sram_2_banks_6_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_2_banks_6_bank_port_1[0] && _zz_sram_2_banks_6_bank_port_2) begin
      sram_2_banks_6_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_6_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_6_bank_port_1[1] && _zz_sram_2_banks_6_bank_port_2) begin
      sram_2_banks_6_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_6_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_6_bank_port_1[2] && _zz_sram_2_banks_6_bank_port_2) begin
      sram_2_banks_6_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_6_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_6_bank_port_1[3] && _zz_sram_2_banks_6_bank_port_2) begin
      sram_2_banks_6_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_6_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_6_banksymbol_read <= sram_2_banks_6_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_6_banksymbol_read_1 <= sram_2_banks_6_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_6_banksymbol_read_2 <= sram_2_banks_6_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_6_banksymbol_read_3 <= sram_2_banks_6_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_7_bank_port1 = {_zz_sram_2_banks_7_banksymbol_read_3, _zz_sram_2_banks_7_banksymbol_read_2, _zz_sram_2_banks_7_banksymbol_read_1, _zz_sram_2_banks_7_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_2_banks_7_bank_port_1[0] && _zz_sram_2_banks_7_bank_port_2) begin
      sram_2_banks_7_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_7_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_7_bank_port_1[1] && _zz_sram_2_banks_7_bank_port_2) begin
      sram_2_banks_7_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_7_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_7_bank_port_1[2] && _zz_sram_2_banks_7_bank_port_2) begin
      sram_2_banks_7_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_7_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_7_bank_port_1[3] && _zz_sram_2_banks_7_bank_port_2) begin
      sram_2_banks_7_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_7_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_7_banksymbol_read <= sram_2_banks_7_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_7_banksymbol_read_1 <= sram_2_banks_7_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_7_banksymbol_read_2 <= sram_2_banks_7_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_7_banksymbol_read_3 <= sram_2_banks_7_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_8_bank_port1 = {_zz_sram_2_banks_8_banksymbol_read_3, _zz_sram_2_banks_8_banksymbol_read_2, _zz_sram_2_banks_8_banksymbol_read_1, _zz_sram_2_banks_8_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_2_banks_8_bank_port_1[0] && _zz_sram_2_banks_8_bank_port_2) begin
      sram_2_banks_8_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_8_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_8_bank_port_1[1] && _zz_sram_2_banks_8_bank_port_2) begin
      sram_2_banks_8_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_8_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_8_bank_port_1[2] && _zz_sram_2_banks_8_bank_port_2) begin
      sram_2_banks_8_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_8_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_8_bank_port_1[3] && _zz_sram_2_banks_8_bank_port_2) begin
      sram_2_banks_8_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_8_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_8_banksymbol_read <= sram_2_banks_8_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_8_banksymbol_read_1 <= sram_2_banks_8_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_8_banksymbol_read_2 <= sram_2_banks_8_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_8_banksymbol_read_3 <= sram_2_banks_8_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_9_bank_port1 = {_zz_sram_2_banks_9_banksymbol_read_3, _zz_sram_2_banks_9_banksymbol_read_2, _zz_sram_2_banks_9_banksymbol_read_1, _zz_sram_2_banks_9_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_2_banks_9_bank_port_1[0] && _zz_sram_2_banks_9_bank_port_2) begin
      sram_2_banks_9_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_9_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_9_bank_port_1[1] && _zz_sram_2_banks_9_bank_port_2) begin
      sram_2_banks_9_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_9_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_9_bank_port_1[2] && _zz_sram_2_banks_9_bank_port_2) begin
      sram_2_banks_9_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_9_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_9_bank_port_1[3] && _zz_sram_2_banks_9_bank_port_2) begin
      sram_2_banks_9_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_9_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_9_banksymbol_read <= sram_2_banks_9_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_9_banksymbol_read_1 <= sram_2_banks_9_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_9_banksymbol_read_2 <= sram_2_banks_9_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_9_banksymbol_read_3 <= sram_2_banks_9_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_10_bank_port1 = {_zz_sram_2_banks_10_banksymbol_read_3, _zz_sram_2_banks_10_banksymbol_read_2, _zz_sram_2_banks_10_banksymbol_read_1, _zz_sram_2_banks_10_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_2_banks_10_bank_port_1[0] && _zz_sram_2_banks_10_bank_port_2) begin
      sram_2_banks_10_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_10_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_10_bank_port_1[1] && _zz_sram_2_banks_10_bank_port_2) begin
      sram_2_banks_10_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_10_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_10_bank_port_1[2] && _zz_sram_2_banks_10_bank_port_2) begin
      sram_2_banks_10_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_10_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_10_bank_port_1[3] && _zz_sram_2_banks_10_bank_port_2) begin
      sram_2_banks_10_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_10_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_10_banksymbol_read <= sram_2_banks_10_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_10_banksymbol_read_1 <= sram_2_banks_10_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_10_banksymbol_read_2 <= sram_2_banks_10_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_10_banksymbol_read_3 <= sram_2_banks_10_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_11_bank_port1 = {_zz_sram_2_banks_11_banksymbol_read_3, _zz_sram_2_banks_11_banksymbol_read_2, _zz_sram_2_banks_11_banksymbol_read_1, _zz_sram_2_banks_11_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_2_banks_11_bank_port_1[0] && _zz_sram_2_banks_11_bank_port_2) begin
      sram_2_banks_11_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_11_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_11_bank_port_1[1] && _zz_sram_2_banks_11_bank_port_2) begin
      sram_2_banks_11_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_11_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_11_bank_port_1[2] && _zz_sram_2_banks_11_bank_port_2) begin
      sram_2_banks_11_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_11_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_11_bank_port_1[3] && _zz_sram_2_banks_11_bank_port_2) begin
      sram_2_banks_11_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_11_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_11_banksymbol_read <= sram_2_banks_11_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_11_banksymbol_read_1 <= sram_2_banks_11_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_11_banksymbol_read_2 <= sram_2_banks_11_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_11_banksymbol_read_3 <= sram_2_banks_11_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_12_bank_port1 = {_zz_sram_2_banks_12_banksymbol_read_3, _zz_sram_2_banks_12_banksymbol_read_2, _zz_sram_2_banks_12_banksymbol_read_1, _zz_sram_2_banks_12_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_2_banks_12_bank_port_1[0] && _zz_sram_2_banks_12_bank_port_2) begin
      sram_2_banks_12_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_12_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_12_bank_port_1[1] && _zz_sram_2_banks_12_bank_port_2) begin
      sram_2_banks_12_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_12_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_12_bank_port_1[2] && _zz_sram_2_banks_12_bank_port_2) begin
      sram_2_banks_12_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_12_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_12_bank_port_1[3] && _zz_sram_2_banks_12_bank_port_2) begin
      sram_2_banks_12_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_12_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_12_banksymbol_read <= sram_2_banks_12_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_12_banksymbol_read_1 <= sram_2_banks_12_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_12_banksymbol_read_2 <= sram_2_banks_12_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_12_banksymbol_read_3 <= sram_2_banks_12_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_13_bank_port1 = {_zz_sram_2_banks_13_banksymbol_read_3, _zz_sram_2_banks_13_banksymbol_read_2, _zz_sram_2_banks_13_banksymbol_read_1, _zz_sram_2_banks_13_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_2_banks_13_bank_port_1[0] && _zz_sram_2_banks_13_bank_port_2) begin
      sram_2_banks_13_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_13_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_13_bank_port_1[1] && _zz_sram_2_banks_13_bank_port_2) begin
      sram_2_banks_13_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_13_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_13_bank_port_1[2] && _zz_sram_2_banks_13_bank_port_2) begin
      sram_2_banks_13_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_13_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_13_bank_port_1[3] && _zz_sram_2_banks_13_bank_port_2) begin
      sram_2_banks_13_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_13_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_13_banksymbol_read <= sram_2_banks_13_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_13_banksymbol_read_1 <= sram_2_banks_13_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_13_banksymbol_read_2 <= sram_2_banks_13_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_13_banksymbol_read_3 <= sram_2_banks_13_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_14_bank_port1 = {_zz_sram_2_banks_14_banksymbol_read_3, _zz_sram_2_banks_14_banksymbol_read_2, _zz_sram_2_banks_14_banksymbol_read_1, _zz_sram_2_banks_14_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_2_banks_14_bank_port_1[0] && _zz_sram_2_banks_14_bank_port_2) begin
      sram_2_banks_14_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_14_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_14_bank_port_1[1] && _zz_sram_2_banks_14_bank_port_2) begin
      sram_2_banks_14_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_14_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_14_bank_port_1[2] && _zz_sram_2_banks_14_bank_port_2) begin
      sram_2_banks_14_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_14_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_14_bank_port_1[3] && _zz_sram_2_banks_14_bank_port_2) begin
      sram_2_banks_14_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_14_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_14_banksymbol_read <= sram_2_banks_14_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_14_banksymbol_read_1 <= sram_2_banks_14_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_14_banksymbol_read_2 <= sram_2_banks_14_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_14_banksymbol_read_3 <= sram_2_banks_14_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_15_bank_port1 = {_zz_sram_2_banks_15_banksymbol_read_3, _zz_sram_2_banks_15_banksymbol_read_2, _zz_sram_2_banks_15_banksymbol_read_1, _zz_sram_2_banks_15_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_2_banks_15_bank_port_1[0] && _zz_sram_2_banks_15_bank_port_2) begin
      sram_2_banks_15_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_15_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_15_bank_port_1[1] && _zz_sram_2_banks_15_bank_port_2) begin
      sram_2_banks_15_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_15_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_15_bank_port_1[2] && _zz_sram_2_banks_15_bank_port_2) begin
      sram_2_banks_15_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_15_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_15_bank_port_1[3] && _zz_sram_2_banks_15_bank_port_2) begin
      sram_2_banks_15_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_15_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_15_banksymbol_read <= sram_2_banks_15_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_15_banksymbol_read_1 <= sram_2_banks_15_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_15_banksymbol_read_2 <= sram_2_banks_15_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_15_banksymbol_read_3 <= sram_2_banks_15_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_0_bank_port1 = {_zz_sram_3_banks_0_banksymbol_read_3, _zz_sram_3_banks_0_banksymbol_read_2, _zz_sram_3_banks_0_banksymbol_read_1, _zz_sram_3_banks_0_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_3_banks_0_bank_port_1[0] && _zz_sram_3_banks_0_bank_port_2) begin
      sram_3_banks_0_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_0_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_0_bank_port_1[1] && _zz_sram_3_banks_0_bank_port_2) begin
      sram_3_banks_0_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_0_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_0_bank_port_1[2] && _zz_sram_3_banks_0_bank_port_2) begin
      sram_3_banks_0_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_0_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_0_bank_port_1[3] && _zz_sram_3_banks_0_bank_port_2) begin
      sram_3_banks_0_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_0_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_0_banksymbol_read <= sram_3_banks_0_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_0_banksymbol_read_1 <= sram_3_banks_0_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_0_banksymbol_read_2 <= sram_3_banks_0_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_0_banksymbol_read_3 <= sram_3_banks_0_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_1_bank_port1 = {_zz_sram_3_banks_1_banksymbol_read_3, _zz_sram_3_banks_1_banksymbol_read_2, _zz_sram_3_banks_1_banksymbol_read_1, _zz_sram_3_banks_1_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_3_banks_1_bank_port_1[0] && _zz_sram_3_banks_1_bank_port_2) begin
      sram_3_banks_1_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_1_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_1_bank_port_1[1] && _zz_sram_3_banks_1_bank_port_2) begin
      sram_3_banks_1_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_1_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_1_bank_port_1[2] && _zz_sram_3_banks_1_bank_port_2) begin
      sram_3_banks_1_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_1_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_1_bank_port_1[3] && _zz_sram_3_banks_1_bank_port_2) begin
      sram_3_banks_1_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_1_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_1_banksymbol_read <= sram_3_banks_1_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_1_banksymbol_read_1 <= sram_3_banks_1_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_1_banksymbol_read_2 <= sram_3_banks_1_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_1_banksymbol_read_3 <= sram_3_banks_1_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_2_bank_port1 = {_zz_sram_3_banks_2_banksymbol_read_3, _zz_sram_3_banks_2_banksymbol_read_2, _zz_sram_3_banks_2_banksymbol_read_1, _zz_sram_3_banks_2_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_3_banks_2_bank_port_1[0] && _zz_sram_3_banks_2_bank_port_2) begin
      sram_3_banks_2_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_2_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_2_bank_port_1[1] && _zz_sram_3_banks_2_bank_port_2) begin
      sram_3_banks_2_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_2_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_2_bank_port_1[2] && _zz_sram_3_banks_2_bank_port_2) begin
      sram_3_banks_2_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_2_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_2_bank_port_1[3] && _zz_sram_3_banks_2_bank_port_2) begin
      sram_3_banks_2_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_2_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_2_banksymbol_read <= sram_3_banks_2_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_2_banksymbol_read_1 <= sram_3_banks_2_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_2_banksymbol_read_2 <= sram_3_banks_2_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_2_banksymbol_read_3 <= sram_3_banks_2_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_3_bank_port1 = {_zz_sram_3_banks_3_banksymbol_read_3, _zz_sram_3_banks_3_banksymbol_read_2, _zz_sram_3_banks_3_banksymbol_read_1, _zz_sram_3_banks_3_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_3_banks_3_bank_port_1[0] && _zz_sram_3_banks_3_bank_port_2) begin
      sram_3_banks_3_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_3_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_3_bank_port_1[1] && _zz_sram_3_banks_3_bank_port_2) begin
      sram_3_banks_3_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_3_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_3_bank_port_1[2] && _zz_sram_3_banks_3_bank_port_2) begin
      sram_3_banks_3_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_3_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_3_bank_port_1[3] && _zz_sram_3_banks_3_bank_port_2) begin
      sram_3_banks_3_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_3_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_3_banksymbol_read <= sram_3_banks_3_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_3_banksymbol_read_1 <= sram_3_banks_3_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_3_banksymbol_read_2 <= sram_3_banks_3_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_3_banksymbol_read_3 <= sram_3_banks_3_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_4_bank_port1 = {_zz_sram_3_banks_4_banksymbol_read_3, _zz_sram_3_banks_4_banksymbol_read_2, _zz_sram_3_banks_4_banksymbol_read_1, _zz_sram_3_banks_4_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_3_banks_4_bank_port_1[0] && _zz_sram_3_banks_4_bank_port_2) begin
      sram_3_banks_4_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_4_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_4_bank_port_1[1] && _zz_sram_3_banks_4_bank_port_2) begin
      sram_3_banks_4_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_4_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_4_bank_port_1[2] && _zz_sram_3_banks_4_bank_port_2) begin
      sram_3_banks_4_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_4_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_4_bank_port_1[3] && _zz_sram_3_banks_4_bank_port_2) begin
      sram_3_banks_4_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_4_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_4_banksymbol_read <= sram_3_banks_4_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_4_banksymbol_read_1 <= sram_3_banks_4_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_4_banksymbol_read_2 <= sram_3_banks_4_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_4_banksymbol_read_3 <= sram_3_banks_4_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_5_bank_port1 = {_zz_sram_3_banks_5_banksymbol_read_3, _zz_sram_3_banks_5_banksymbol_read_2, _zz_sram_3_banks_5_banksymbol_read_1, _zz_sram_3_banks_5_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_3_banks_5_bank_port_1[0] && _zz_sram_3_banks_5_bank_port_2) begin
      sram_3_banks_5_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_5_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_5_bank_port_1[1] && _zz_sram_3_banks_5_bank_port_2) begin
      sram_3_banks_5_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_5_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_5_bank_port_1[2] && _zz_sram_3_banks_5_bank_port_2) begin
      sram_3_banks_5_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_5_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_5_bank_port_1[3] && _zz_sram_3_banks_5_bank_port_2) begin
      sram_3_banks_5_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_5_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_5_banksymbol_read <= sram_3_banks_5_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_5_banksymbol_read_1 <= sram_3_banks_5_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_5_banksymbol_read_2 <= sram_3_banks_5_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_5_banksymbol_read_3 <= sram_3_banks_5_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_6_bank_port1 = {_zz_sram_3_banks_6_banksymbol_read_3, _zz_sram_3_banks_6_banksymbol_read_2, _zz_sram_3_banks_6_banksymbol_read_1, _zz_sram_3_banks_6_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_3_banks_6_bank_port_1[0] && _zz_sram_3_banks_6_bank_port_2) begin
      sram_3_banks_6_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_6_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_6_bank_port_1[1] && _zz_sram_3_banks_6_bank_port_2) begin
      sram_3_banks_6_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_6_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_6_bank_port_1[2] && _zz_sram_3_banks_6_bank_port_2) begin
      sram_3_banks_6_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_6_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_6_bank_port_1[3] && _zz_sram_3_banks_6_bank_port_2) begin
      sram_3_banks_6_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_6_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_6_banksymbol_read <= sram_3_banks_6_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_6_banksymbol_read_1 <= sram_3_banks_6_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_6_banksymbol_read_2 <= sram_3_banks_6_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_6_banksymbol_read_3 <= sram_3_banks_6_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_7_bank_port1 = {_zz_sram_3_banks_7_banksymbol_read_3, _zz_sram_3_banks_7_banksymbol_read_2, _zz_sram_3_banks_7_banksymbol_read_1, _zz_sram_3_banks_7_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_3_banks_7_bank_port_1[0] && _zz_sram_3_banks_7_bank_port_2) begin
      sram_3_banks_7_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_7_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_7_bank_port_1[1] && _zz_sram_3_banks_7_bank_port_2) begin
      sram_3_banks_7_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_7_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_7_bank_port_1[2] && _zz_sram_3_banks_7_bank_port_2) begin
      sram_3_banks_7_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_7_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_7_bank_port_1[3] && _zz_sram_3_banks_7_bank_port_2) begin
      sram_3_banks_7_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_7_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_7_banksymbol_read <= sram_3_banks_7_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_7_banksymbol_read_1 <= sram_3_banks_7_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_7_banksymbol_read_2 <= sram_3_banks_7_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_7_banksymbol_read_3 <= sram_3_banks_7_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_8_bank_port1 = {_zz_sram_3_banks_8_banksymbol_read_3, _zz_sram_3_banks_8_banksymbol_read_2, _zz_sram_3_banks_8_banksymbol_read_1, _zz_sram_3_banks_8_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_3_banks_8_bank_port_1[0] && _zz_sram_3_banks_8_bank_port_2) begin
      sram_3_banks_8_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_8_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_8_bank_port_1[1] && _zz_sram_3_banks_8_bank_port_2) begin
      sram_3_banks_8_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_8_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_8_bank_port_1[2] && _zz_sram_3_banks_8_bank_port_2) begin
      sram_3_banks_8_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_8_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_8_bank_port_1[3] && _zz_sram_3_banks_8_bank_port_2) begin
      sram_3_banks_8_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_8_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_8_banksymbol_read <= sram_3_banks_8_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_8_banksymbol_read_1 <= sram_3_banks_8_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_8_banksymbol_read_2 <= sram_3_banks_8_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_8_banksymbol_read_3 <= sram_3_banks_8_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_9_bank_port1 = {_zz_sram_3_banks_9_banksymbol_read_3, _zz_sram_3_banks_9_banksymbol_read_2, _zz_sram_3_banks_9_banksymbol_read_1, _zz_sram_3_banks_9_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_3_banks_9_bank_port_1[0] && _zz_sram_3_banks_9_bank_port_2) begin
      sram_3_banks_9_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_9_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_9_bank_port_1[1] && _zz_sram_3_banks_9_bank_port_2) begin
      sram_3_banks_9_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_9_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_9_bank_port_1[2] && _zz_sram_3_banks_9_bank_port_2) begin
      sram_3_banks_9_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_9_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_9_bank_port_1[3] && _zz_sram_3_banks_9_bank_port_2) begin
      sram_3_banks_9_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_9_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_9_banksymbol_read <= sram_3_banks_9_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_9_banksymbol_read_1 <= sram_3_banks_9_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_9_banksymbol_read_2 <= sram_3_banks_9_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_9_banksymbol_read_3 <= sram_3_banks_9_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_10_bank_port1 = {_zz_sram_3_banks_10_banksymbol_read_3, _zz_sram_3_banks_10_banksymbol_read_2, _zz_sram_3_banks_10_banksymbol_read_1, _zz_sram_3_banks_10_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_3_banks_10_bank_port_1[0] && _zz_sram_3_banks_10_bank_port_2) begin
      sram_3_banks_10_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_10_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_10_bank_port_1[1] && _zz_sram_3_banks_10_bank_port_2) begin
      sram_3_banks_10_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_10_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_10_bank_port_1[2] && _zz_sram_3_banks_10_bank_port_2) begin
      sram_3_banks_10_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_10_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_10_bank_port_1[3] && _zz_sram_3_banks_10_bank_port_2) begin
      sram_3_banks_10_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_10_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_10_banksymbol_read <= sram_3_banks_10_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_10_banksymbol_read_1 <= sram_3_banks_10_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_10_banksymbol_read_2 <= sram_3_banks_10_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_10_banksymbol_read_3 <= sram_3_banks_10_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_11_bank_port1 = {_zz_sram_3_banks_11_banksymbol_read_3, _zz_sram_3_banks_11_banksymbol_read_2, _zz_sram_3_banks_11_banksymbol_read_1, _zz_sram_3_banks_11_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_3_banks_11_bank_port_1[0] && _zz_sram_3_banks_11_bank_port_2) begin
      sram_3_banks_11_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_11_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_11_bank_port_1[1] && _zz_sram_3_banks_11_bank_port_2) begin
      sram_3_banks_11_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_11_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_11_bank_port_1[2] && _zz_sram_3_banks_11_bank_port_2) begin
      sram_3_banks_11_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_11_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_11_bank_port_1[3] && _zz_sram_3_banks_11_bank_port_2) begin
      sram_3_banks_11_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_11_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_11_banksymbol_read <= sram_3_banks_11_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_11_banksymbol_read_1 <= sram_3_banks_11_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_11_banksymbol_read_2 <= sram_3_banks_11_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_11_banksymbol_read_3 <= sram_3_banks_11_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_12_bank_port1 = {_zz_sram_3_banks_12_banksymbol_read_3, _zz_sram_3_banks_12_banksymbol_read_2, _zz_sram_3_banks_12_banksymbol_read_1, _zz_sram_3_banks_12_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_3_banks_12_bank_port_1[0] && _zz_sram_3_banks_12_bank_port_2) begin
      sram_3_banks_12_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_12_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_12_bank_port_1[1] && _zz_sram_3_banks_12_bank_port_2) begin
      sram_3_banks_12_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_12_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_12_bank_port_1[2] && _zz_sram_3_banks_12_bank_port_2) begin
      sram_3_banks_12_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_12_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_12_bank_port_1[3] && _zz_sram_3_banks_12_bank_port_2) begin
      sram_3_banks_12_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_12_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_12_banksymbol_read <= sram_3_banks_12_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_12_banksymbol_read_1 <= sram_3_banks_12_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_12_banksymbol_read_2 <= sram_3_banks_12_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_12_banksymbol_read_3 <= sram_3_banks_12_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_13_bank_port1 = {_zz_sram_3_banks_13_banksymbol_read_3, _zz_sram_3_banks_13_banksymbol_read_2, _zz_sram_3_banks_13_banksymbol_read_1, _zz_sram_3_banks_13_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_3_banks_13_bank_port_1[0] && _zz_sram_3_banks_13_bank_port_2) begin
      sram_3_banks_13_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_13_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_13_bank_port_1[1] && _zz_sram_3_banks_13_bank_port_2) begin
      sram_3_banks_13_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_13_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_13_bank_port_1[2] && _zz_sram_3_banks_13_bank_port_2) begin
      sram_3_banks_13_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_13_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_13_bank_port_1[3] && _zz_sram_3_banks_13_bank_port_2) begin
      sram_3_banks_13_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_13_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_13_banksymbol_read <= sram_3_banks_13_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_13_banksymbol_read_1 <= sram_3_banks_13_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_13_banksymbol_read_2 <= sram_3_banks_13_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_13_banksymbol_read_3 <= sram_3_banks_13_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_14_bank_port1 = {_zz_sram_3_banks_14_banksymbol_read_3, _zz_sram_3_banks_14_banksymbol_read_2, _zz_sram_3_banks_14_banksymbol_read_1, _zz_sram_3_banks_14_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_3_banks_14_bank_port_1[0] && _zz_sram_3_banks_14_bank_port_2) begin
      sram_3_banks_14_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_14_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_14_bank_port_1[1] && _zz_sram_3_banks_14_bank_port_2) begin
      sram_3_banks_14_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_14_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_14_bank_port_1[2] && _zz_sram_3_banks_14_bank_port_2) begin
      sram_3_banks_14_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_14_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_14_bank_port_1[3] && _zz_sram_3_banks_14_bank_port_2) begin
      sram_3_banks_14_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_14_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_14_banksymbol_read <= sram_3_banks_14_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_14_banksymbol_read_1 <= sram_3_banks_14_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_14_banksymbol_read_2 <= sram_3_banks_14_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_14_banksymbol_read_3 <= sram_3_banks_14_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_15_bank_port1 = {_zz_sram_3_banks_15_banksymbol_read_3, _zz_sram_3_banks_15_banksymbol_read_2, _zz_sram_3_banks_15_banksymbol_read_1, _zz_sram_3_banks_15_banksymbol_read};
  end
  always @(posedge io_axiClk) begin
    if(_zz_sram_3_banks_15_bank_port_1[0] && _zz_sram_3_banks_15_bank_port_2) begin
      sram_3_banks_15_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_15_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_15_bank_port_1[1] && _zz_sram_3_banks_15_bank_port_2) begin
      sram_3_banks_15_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_15_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_15_bank_port_1[2] && _zz_sram_3_banks_15_bank_port_2) begin
      sram_3_banks_15_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_15_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_15_bank_port_1[3] && _zz_sram_3_banks_15_bank_port_2) begin
      sram_3_banks_15_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_15_bank_port[31 : 24];
    end
  end

  always @(posedge io_axiClk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_15_banksymbol_read <= sram_3_banks_15_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_15_banksymbol_read_1 <= sram_3_banks_15_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_15_banksymbol_read_2 <= sram_3_banks_15_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_15_banksymbol_read_3 <= sram_3_banks_15_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    sram_0_ports_rsp_payload_data[31 : 0] = _zz_sram_0_banks_0_bank_port1;
    sram_0_ports_rsp_payload_data[63 : 32] = _zz_sram_0_banks_1_bank_port1;
    sram_0_ports_rsp_payload_data[95 : 64] = _zz_sram_0_banks_2_bank_port1;
    sram_0_ports_rsp_payload_data[127 : 96] = _zz_sram_0_banks_3_bank_port1;
    sram_0_ports_rsp_payload_data[159 : 128] = _zz_sram_0_banks_4_bank_port1;
    sram_0_ports_rsp_payload_data[191 : 160] = _zz_sram_0_banks_5_bank_port1;
    sram_0_ports_rsp_payload_data[223 : 192] = _zz_sram_0_banks_6_bank_port1;
    sram_0_ports_rsp_payload_data[255 : 224] = _zz_sram_0_banks_7_bank_port1;
    sram_0_ports_rsp_payload_data[287 : 256] = _zz_sram_0_banks_8_bank_port1;
    sram_0_ports_rsp_payload_data[319 : 288] = _zz_sram_0_banks_9_bank_port1;
    sram_0_ports_rsp_payload_data[351 : 320] = _zz_sram_0_banks_10_bank_port1;
    sram_0_ports_rsp_payload_data[383 : 352] = _zz_sram_0_banks_11_bank_port1;
    sram_0_ports_rsp_payload_data[415 : 384] = _zz_sram_0_banks_12_bank_port1;
    sram_0_ports_rsp_payload_data[447 : 416] = _zz_sram_0_banks_13_bank_port1;
    sram_0_ports_rsp_payload_data[479 : 448] = _zz_sram_0_banks_14_bank_port1;
    sram_0_ports_rsp_payload_data[511 : 480] = _zz_sram_0_banks_15_bank_port1;
  end

  assign when_SramBanks_l66 = (sram_0_ports_cmd_valid && (sram_0_ports_cmd_payload_wen == 16'h0));
  assign sram_0_ports_rsp_valid = _zz_sram_0_ports_rsp_valid;
  always @(*) begin
    sram_1_ports_rsp_payload_data[31 : 0] = _zz_sram_1_banks_0_bank_port1;
    sram_1_ports_rsp_payload_data[63 : 32] = _zz_sram_1_banks_1_bank_port1;
    sram_1_ports_rsp_payload_data[95 : 64] = _zz_sram_1_banks_2_bank_port1;
    sram_1_ports_rsp_payload_data[127 : 96] = _zz_sram_1_banks_3_bank_port1;
    sram_1_ports_rsp_payload_data[159 : 128] = _zz_sram_1_banks_4_bank_port1;
    sram_1_ports_rsp_payload_data[191 : 160] = _zz_sram_1_banks_5_bank_port1;
    sram_1_ports_rsp_payload_data[223 : 192] = _zz_sram_1_banks_6_bank_port1;
    sram_1_ports_rsp_payload_data[255 : 224] = _zz_sram_1_banks_7_bank_port1;
    sram_1_ports_rsp_payload_data[287 : 256] = _zz_sram_1_banks_8_bank_port1;
    sram_1_ports_rsp_payload_data[319 : 288] = _zz_sram_1_banks_9_bank_port1;
    sram_1_ports_rsp_payload_data[351 : 320] = _zz_sram_1_banks_10_bank_port1;
    sram_1_ports_rsp_payload_data[383 : 352] = _zz_sram_1_banks_11_bank_port1;
    sram_1_ports_rsp_payload_data[415 : 384] = _zz_sram_1_banks_12_bank_port1;
    sram_1_ports_rsp_payload_data[447 : 416] = _zz_sram_1_banks_13_bank_port1;
    sram_1_ports_rsp_payload_data[479 : 448] = _zz_sram_1_banks_14_bank_port1;
    sram_1_ports_rsp_payload_data[511 : 480] = _zz_sram_1_banks_15_bank_port1;
  end

  assign when_SramBanks_l66_1 = (sram_1_ports_cmd_valid && (sram_1_ports_cmd_payload_wen == 16'h0));
  assign sram_1_ports_rsp_valid = _zz_sram_1_ports_rsp_valid;
  always @(*) begin
    sram_2_ports_rsp_payload_data[31 : 0] = _zz_sram_2_banks_0_bank_port1;
    sram_2_ports_rsp_payload_data[63 : 32] = _zz_sram_2_banks_1_bank_port1;
    sram_2_ports_rsp_payload_data[95 : 64] = _zz_sram_2_banks_2_bank_port1;
    sram_2_ports_rsp_payload_data[127 : 96] = _zz_sram_2_banks_3_bank_port1;
    sram_2_ports_rsp_payload_data[159 : 128] = _zz_sram_2_banks_4_bank_port1;
    sram_2_ports_rsp_payload_data[191 : 160] = _zz_sram_2_banks_5_bank_port1;
    sram_2_ports_rsp_payload_data[223 : 192] = _zz_sram_2_banks_6_bank_port1;
    sram_2_ports_rsp_payload_data[255 : 224] = _zz_sram_2_banks_7_bank_port1;
    sram_2_ports_rsp_payload_data[287 : 256] = _zz_sram_2_banks_8_bank_port1;
    sram_2_ports_rsp_payload_data[319 : 288] = _zz_sram_2_banks_9_bank_port1;
    sram_2_ports_rsp_payload_data[351 : 320] = _zz_sram_2_banks_10_bank_port1;
    sram_2_ports_rsp_payload_data[383 : 352] = _zz_sram_2_banks_11_bank_port1;
    sram_2_ports_rsp_payload_data[415 : 384] = _zz_sram_2_banks_12_bank_port1;
    sram_2_ports_rsp_payload_data[447 : 416] = _zz_sram_2_banks_13_bank_port1;
    sram_2_ports_rsp_payload_data[479 : 448] = _zz_sram_2_banks_14_bank_port1;
    sram_2_ports_rsp_payload_data[511 : 480] = _zz_sram_2_banks_15_bank_port1;
  end

  assign when_SramBanks_l66_2 = (sram_2_ports_cmd_valid && (sram_2_ports_cmd_payload_wen == 16'h0));
  assign sram_2_ports_rsp_valid = _zz_sram_2_ports_rsp_valid;
  always @(*) begin
    sram_3_ports_rsp_payload_data[31 : 0] = _zz_sram_3_banks_0_bank_port1;
    sram_3_ports_rsp_payload_data[63 : 32] = _zz_sram_3_banks_1_bank_port1;
    sram_3_ports_rsp_payload_data[95 : 64] = _zz_sram_3_banks_2_bank_port1;
    sram_3_ports_rsp_payload_data[127 : 96] = _zz_sram_3_banks_3_bank_port1;
    sram_3_ports_rsp_payload_data[159 : 128] = _zz_sram_3_banks_4_bank_port1;
    sram_3_ports_rsp_payload_data[191 : 160] = _zz_sram_3_banks_5_bank_port1;
    sram_3_ports_rsp_payload_data[223 : 192] = _zz_sram_3_banks_6_bank_port1;
    sram_3_ports_rsp_payload_data[255 : 224] = _zz_sram_3_banks_7_bank_port1;
    sram_3_ports_rsp_payload_data[287 : 256] = _zz_sram_3_banks_8_bank_port1;
    sram_3_ports_rsp_payload_data[319 : 288] = _zz_sram_3_banks_9_bank_port1;
    sram_3_ports_rsp_payload_data[351 : 320] = _zz_sram_3_banks_10_bank_port1;
    sram_3_ports_rsp_payload_data[383 : 352] = _zz_sram_3_banks_11_bank_port1;
    sram_3_ports_rsp_payload_data[415 : 384] = _zz_sram_3_banks_12_bank_port1;
    sram_3_ports_rsp_payload_data[447 : 416] = _zz_sram_3_banks_13_bank_port1;
    sram_3_ports_rsp_payload_data[479 : 448] = _zz_sram_3_banks_14_bank_port1;
    sram_3_ports_rsp_payload_data[511 : 480] = _zz_sram_3_banks_15_bank_port1;
  end

  assign when_SramBanks_l66_3 = (sram_3_ports_cmd_valid && (sram_3_ports_cmd_payload_wen == 16'h0));
  assign sram_3_ports_rsp_valid = _zz_sram_3_ports_rsp_valid;
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      _zz_sram_0_ports_rsp_valid <= 1'b0;
      _zz_sram_1_ports_rsp_valid <= 1'b0;
      _zz_sram_2_ports_rsp_valid <= 1'b0;
      _zz_sram_3_ports_rsp_valid <= 1'b0;
    end else begin
      if(when_SramBanks_l66) begin
        _zz_sram_0_ports_rsp_valid <= 1'b1;
      end else begin
        _zz_sram_0_ports_rsp_valid <= 1'b0;
      end
      if(when_SramBanks_l66_1) begin
        _zz_sram_1_ports_rsp_valid <= 1'b1;
      end else begin
        _zz_sram_1_ports_rsp_valid <= 1'b0;
      end
      if(when_SramBanks_l66_2) begin
        _zz_sram_2_ports_rsp_valid <= 1'b1;
      end else begin
        _zz_sram_2_ports_rsp_valid <= 1'b0;
      end
      if(when_SramBanks_l66_3) begin
        _zz_sram_3_ports_rsp_valid <= 1'b1;
      end else begin
        _zz_sram_3_ports_rsp_valid <= 1'b0;
      end
    end
  end


endmodule

module ICache (
  input               flush,
  input               cpu_cmd_valid,
  output              cpu_cmd_ready,
  input      [63:0]   cpu_cmd_payload_addr,
  output              cpu_rsp_valid,
  output     [31:0]   cpu_rsp_payload_data,
  output reg          sram_0_ports_cmd_valid,
  output reg [3:0]    sram_0_ports_cmd_payload_addr,
  output reg [15:0]   sram_0_ports_cmd_payload_wen,
  output reg [511:0]  sram_0_ports_cmd_payload_wdata,
  output reg [63:0]   sram_0_ports_cmd_payload_wstrb,
  input               sram_0_ports_rsp_valid,
  input      [511:0]  sram_0_ports_rsp_payload_data,
  output reg          sram_1_ports_cmd_valid,
  output reg [3:0]    sram_1_ports_cmd_payload_addr,
  output reg [15:0]   sram_1_ports_cmd_payload_wen,
  output reg [511:0]  sram_1_ports_cmd_payload_wdata,
  output reg [63:0]   sram_1_ports_cmd_payload_wstrb,
  input               sram_1_ports_rsp_valid,
  input      [511:0]  sram_1_ports_rsp_payload_data,
  output reg          sram_2_ports_cmd_valid,
  output reg [3:0]    sram_2_ports_cmd_payload_addr,
  output reg [15:0]   sram_2_ports_cmd_payload_wen,
  output reg [511:0]  sram_2_ports_cmd_payload_wdata,
  output reg [63:0]   sram_2_ports_cmd_payload_wstrb,
  input               sram_2_ports_rsp_valid,
  input      [511:0]  sram_2_ports_rsp_payload_data,
  output reg          sram_3_ports_cmd_valid,
  output reg [3:0]    sram_3_ports_cmd_payload_addr,
  output reg [15:0]   sram_3_ports_cmd_payload_wen,
  output reg [511:0]  sram_3_ports_cmd_payload_wdata,
  output reg [63:0]   sram_3_ports_cmd_payload_wstrb,
  input               sram_3_ports_rsp_valid,
  input      [511:0]  sram_3_ports_rsp_payload_data,
  output              next_level_cmd_valid,
  input               next_level_cmd_ready,
  output     [63:0]   next_level_cmd_payload_addr,
  output     [3:0]    next_level_cmd_payload_len,
  output     [2:0]    next_level_cmd_payload_size,
  input               next_level_rsp_valid,
  input      [63:0]   next_level_rsp_payload_data,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  wire       [3:0]    _zz_flush_cnt_valueNext;
  wire       [0:0]    _zz_flush_cnt_valueNext_1;
  wire       [2:0]    _zz_next_level_data_cnt_valueNext;
  wire       [0:0]    _zz_next_level_data_cnt_valueNext_1;
  wire       [7:0]    _zz__zz_cache_hit_gnt_0_3;
  wire       [7:0]    _zz__zz_cache_hit_gnt_0_3_1;
  wire       [3:0]    _zz__zz_cache_hit_gnt_0_3_2;
  wire       [7:0]    _zz__zz_cache_invld_gnt_0_3;
  wire       [7:0]    _zz__zz_cache_invld_gnt_0_3_1;
  wire       [3:0]    _zz__zz_cache_invld_gnt_0_3_2;
  wire       [7:0]    _zz__zz_cache_victim_gnt_0_3;
  wire       [7:0]    _zz__zz_cache_victim_gnt_0_3_1;
  wire       [3:0]    _zz__zz_cache_victim_gnt_0_3_2;
  reg        [53:0]   _zz_cache_tag_0;
  reg                 _zz_cache_hit_0;
  reg                 _zz_cache_mru_0;
  reg                 _zz_cache_invld_d1_0;
  reg                 _zz_cache_lru_d1_0;
  wire       [4:0]    _zz_sram_0_ports_cmd_payload_wen_1;
  wire       [9:0]    _zz_sram_0_ports_cmd_payload_wdata;
  wire       [9:0]    _zz_sram_0_ports_cmd_payload_wstrb;
  wire       [9:0]    _zz_sram_0_ports_cmd_payload_wstrb_1;
  reg        [53:0]   _zz_cache_tag_1;
  reg                 _zz_cache_hit_1;
  reg                 _zz_cache_mru_1;
  reg                 _zz_cache_invld_d1_1;
  reg                 _zz_cache_lru_d1_1;
  wire       [4:0]    _zz_sram_1_ports_cmd_payload_wen_1;
  wire       [9:0]    _zz_sram_1_ports_cmd_payload_wdata;
  wire       [9:0]    _zz_sram_1_ports_cmd_payload_wstrb;
  wire       [9:0]    _zz_sram_1_ports_cmd_payload_wstrb_1;
  reg        [53:0]   _zz_cache_tag_2;
  reg                 _zz_cache_hit_2;
  reg                 _zz_cache_mru_2;
  reg                 _zz_cache_invld_d1_2;
  reg                 _zz_cache_lru_d1_2;
  wire       [4:0]    _zz_sram_2_ports_cmd_payload_wen_1;
  wire       [9:0]    _zz_sram_2_ports_cmd_payload_wdata;
  wire       [9:0]    _zz_sram_2_ports_cmd_payload_wstrb;
  wire       [9:0]    _zz_sram_2_ports_cmd_payload_wstrb_1;
  reg        [53:0]   _zz_cache_tag_3;
  reg                 _zz_cache_hit_3;
  reg                 _zz_cache_mru_3;
  reg                 _zz_cache_invld_d1_3;
  reg                 _zz_cache_lru_d1_3;
  wire       [4:0]    _zz_sram_3_ports_cmd_payload_wen_1;
  wire       [9:0]    _zz_sram_3_ports_cmd_payload_wdata;
  wire       [9:0]    _zz_sram_3_ports_cmd_payload_wstrb;
  wire       [9:0]    _zz_sram_3_ports_cmd_payload_wstrb_1;
  reg        [511:0]  _zz__zz_hit_data;
  reg        [31:0]   _zz_hit_data_1;
  reg        [511:0]  _zz__zz_miss_data;
  reg        [31:0]   _zz_miss_data_1;
  reg                 _zz_cpu_rsp_valid;
  reg                 _zz_cpu_rsp_valid_1;
  reg                 ways_0_metas_0_vld;
  reg        [53:0]   ways_0_metas_0_tag;
  reg                 ways_0_metas_0_mru;
  reg                 ways_0_metas_1_vld;
  reg        [53:0]   ways_0_metas_1_tag;
  reg                 ways_0_metas_1_mru;
  reg                 ways_0_metas_2_vld;
  reg        [53:0]   ways_0_metas_2_tag;
  reg                 ways_0_metas_2_mru;
  reg                 ways_0_metas_3_vld;
  reg        [53:0]   ways_0_metas_3_tag;
  reg                 ways_0_metas_3_mru;
  reg                 ways_0_metas_4_vld;
  reg        [53:0]   ways_0_metas_4_tag;
  reg                 ways_0_metas_4_mru;
  reg                 ways_0_metas_5_vld;
  reg        [53:0]   ways_0_metas_5_tag;
  reg                 ways_0_metas_5_mru;
  reg                 ways_0_metas_6_vld;
  reg        [53:0]   ways_0_metas_6_tag;
  reg                 ways_0_metas_6_mru;
  reg                 ways_0_metas_7_vld;
  reg        [53:0]   ways_0_metas_7_tag;
  reg                 ways_0_metas_7_mru;
  reg                 ways_0_metas_8_vld;
  reg        [53:0]   ways_0_metas_8_tag;
  reg                 ways_0_metas_8_mru;
  reg                 ways_0_metas_9_vld;
  reg        [53:0]   ways_0_metas_9_tag;
  reg                 ways_0_metas_9_mru;
  reg                 ways_0_metas_10_vld;
  reg        [53:0]   ways_0_metas_10_tag;
  reg                 ways_0_metas_10_mru;
  reg                 ways_0_metas_11_vld;
  reg        [53:0]   ways_0_metas_11_tag;
  reg                 ways_0_metas_11_mru;
  reg                 ways_0_metas_12_vld;
  reg        [53:0]   ways_0_metas_12_tag;
  reg                 ways_0_metas_12_mru;
  reg                 ways_0_metas_13_vld;
  reg        [53:0]   ways_0_metas_13_tag;
  reg                 ways_0_metas_13_mru;
  reg                 ways_0_metas_14_vld;
  reg        [53:0]   ways_0_metas_14_tag;
  reg                 ways_0_metas_14_mru;
  reg                 ways_0_metas_15_vld;
  reg        [53:0]   ways_0_metas_15_tag;
  reg                 ways_0_metas_15_mru;
  reg                 ways_1_metas_0_vld;
  reg        [53:0]   ways_1_metas_0_tag;
  reg                 ways_1_metas_0_mru;
  reg                 ways_1_metas_1_vld;
  reg        [53:0]   ways_1_metas_1_tag;
  reg                 ways_1_metas_1_mru;
  reg                 ways_1_metas_2_vld;
  reg        [53:0]   ways_1_metas_2_tag;
  reg                 ways_1_metas_2_mru;
  reg                 ways_1_metas_3_vld;
  reg        [53:0]   ways_1_metas_3_tag;
  reg                 ways_1_metas_3_mru;
  reg                 ways_1_metas_4_vld;
  reg        [53:0]   ways_1_metas_4_tag;
  reg                 ways_1_metas_4_mru;
  reg                 ways_1_metas_5_vld;
  reg        [53:0]   ways_1_metas_5_tag;
  reg                 ways_1_metas_5_mru;
  reg                 ways_1_metas_6_vld;
  reg        [53:0]   ways_1_metas_6_tag;
  reg                 ways_1_metas_6_mru;
  reg                 ways_1_metas_7_vld;
  reg        [53:0]   ways_1_metas_7_tag;
  reg                 ways_1_metas_7_mru;
  reg                 ways_1_metas_8_vld;
  reg        [53:0]   ways_1_metas_8_tag;
  reg                 ways_1_metas_8_mru;
  reg                 ways_1_metas_9_vld;
  reg        [53:0]   ways_1_metas_9_tag;
  reg                 ways_1_metas_9_mru;
  reg                 ways_1_metas_10_vld;
  reg        [53:0]   ways_1_metas_10_tag;
  reg                 ways_1_metas_10_mru;
  reg                 ways_1_metas_11_vld;
  reg        [53:0]   ways_1_metas_11_tag;
  reg                 ways_1_metas_11_mru;
  reg                 ways_1_metas_12_vld;
  reg        [53:0]   ways_1_metas_12_tag;
  reg                 ways_1_metas_12_mru;
  reg                 ways_1_metas_13_vld;
  reg        [53:0]   ways_1_metas_13_tag;
  reg                 ways_1_metas_13_mru;
  reg                 ways_1_metas_14_vld;
  reg        [53:0]   ways_1_metas_14_tag;
  reg                 ways_1_metas_14_mru;
  reg                 ways_1_metas_15_vld;
  reg        [53:0]   ways_1_metas_15_tag;
  reg                 ways_1_metas_15_mru;
  reg                 ways_2_metas_0_vld;
  reg        [53:0]   ways_2_metas_0_tag;
  reg                 ways_2_metas_0_mru;
  reg                 ways_2_metas_1_vld;
  reg        [53:0]   ways_2_metas_1_tag;
  reg                 ways_2_metas_1_mru;
  reg                 ways_2_metas_2_vld;
  reg        [53:0]   ways_2_metas_2_tag;
  reg                 ways_2_metas_2_mru;
  reg                 ways_2_metas_3_vld;
  reg        [53:0]   ways_2_metas_3_tag;
  reg                 ways_2_metas_3_mru;
  reg                 ways_2_metas_4_vld;
  reg        [53:0]   ways_2_metas_4_tag;
  reg                 ways_2_metas_4_mru;
  reg                 ways_2_metas_5_vld;
  reg        [53:0]   ways_2_metas_5_tag;
  reg                 ways_2_metas_5_mru;
  reg                 ways_2_metas_6_vld;
  reg        [53:0]   ways_2_metas_6_tag;
  reg                 ways_2_metas_6_mru;
  reg                 ways_2_metas_7_vld;
  reg        [53:0]   ways_2_metas_7_tag;
  reg                 ways_2_metas_7_mru;
  reg                 ways_2_metas_8_vld;
  reg        [53:0]   ways_2_metas_8_tag;
  reg                 ways_2_metas_8_mru;
  reg                 ways_2_metas_9_vld;
  reg        [53:0]   ways_2_metas_9_tag;
  reg                 ways_2_metas_9_mru;
  reg                 ways_2_metas_10_vld;
  reg        [53:0]   ways_2_metas_10_tag;
  reg                 ways_2_metas_10_mru;
  reg                 ways_2_metas_11_vld;
  reg        [53:0]   ways_2_metas_11_tag;
  reg                 ways_2_metas_11_mru;
  reg                 ways_2_metas_12_vld;
  reg        [53:0]   ways_2_metas_12_tag;
  reg                 ways_2_metas_12_mru;
  reg                 ways_2_metas_13_vld;
  reg        [53:0]   ways_2_metas_13_tag;
  reg                 ways_2_metas_13_mru;
  reg                 ways_2_metas_14_vld;
  reg        [53:0]   ways_2_metas_14_tag;
  reg                 ways_2_metas_14_mru;
  reg                 ways_2_metas_15_vld;
  reg        [53:0]   ways_2_metas_15_tag;
  reg                 ways_2_metas_15_mru;
  reg                 ways_3_metas_0_vld;
  reg        [53:0]   ways_3_metas_0_tag;
  reg                 ways_3_metas_0_mru;
  reg                 ways_3_metas_1_vld;
  reg        [53:0]   ways_3_metas_1_tag;
  reg                 ways_3_metas_1_mru;
  reg                 ways_3_metas_2_vld;
  reg        [53:0]   ways_3_metas_2_tag;
  reg                 ways_3_metas_2_mru;
  reg                 ways_3_metas_3_vld;
  reg        [53:0]   ways_3_metas_3_tag;
  reg                 ways_3_metas_3_mru;
  reg                 ways_3_metas_4_vld;
  reg        [53:0]   ways_3_metas_4_tag;
  reg                 ways_3_metas_4_mru;
  reg                 ways_3_metas_5_vld;
  reg        [53:0]   ways_3_metas_5_tag;
  reg                 ways_3_metas_5_mru;
  reg                 ways_3_metas_6_vld;
  reg        [53:0]   ways_3_metas_6_tag;
  reg                 ways_3_metas_6_mru;
  reg                 ways_3_metas_7_vld;
  reg        [53:0]   ways_3_metas_7_tag;
  reg                 ways_3_metas_7_mru;
  reg                 ways_3_metas_8_vld;
  reg        [53:0]   ways_3_metas_8_tag;
  reg                 ways_3_metas_8_mru;
  reg                 ways_3_metas_9_vld;
  reg        [53:0]   ways_3_metas_9_tag;
  reg                 ways_3_metas_9_mru;
  reg                 ways_3_metas_10_vld;
  reg        [53:0]   ways_3_metas_10_tag;
  reg                 ways_3_metas_10_mru;
  reg                 ways_3_metas_11_vld;
  reg        [53:0]   ways_3_metas_11_tag;
  reg                 ways_3_metas_11_mru;
  reg                 ways_3_metas_12_vld;
  reg        [53:0]   ways_3_metas_12_tag;
  reg                 ways_3_metas_12_mru;
  reg                 ways_3_metas_13_vld;
  reg        [53:0]   ways_3_metas_13_tag;
  reg                 ways_3_metas_13_mru;
  reg                 ways_3_metas_14_vld;
  reg        [53:0]   ways_3_metas_14_tag;
  reg                 ways_3_metas_14_mru;
  reg                 ways_3_metas_15_vld;
  reg        [53:0]   ways_3_metas_15_tag;
  reg                 ways_3_metas_15_mru;
  wire       [53:0]   cache_tag_0;
  wire       [53:0]   cache_tag_1;
  wire       [53:0]   cache_tag_2;
  wire       [53:0]   cache_tag_3;
  wire                cache_hit_0;
  wire                cache_hit_1;
  wire                cache_hit_2;
  wire                cache_hit_3;
  wire                cache_invld_d1_0;
  wire                cache_invld_d1_1;
  wire                cache_invld_d1_2;
  wire                cache_invld_d1_3;
  wire                cache_victim_0;
  wire                cache_victim_1;
  wire                cache_victim_2;
  wire                cache_victim_3;
  wire                cache_mru_0;
  wire                cache_mru_1;
  wire                cache_mru_2;
  wire                cache_mru_3;
  wire                cache_lru_d1_0;
  wire                cache_lru_d1_1;
  wire                cache_lru_d1_2;
  wire                cache_lru_d1_3;
  wire       [1:0]    hit_id;
  reg        [1:0]    hit_id_d1;
  wire       [1:0]    evict_id;
  wire       [1:0]    invld_id;
  wire       [1:0]    victim_id;
  wire                mru_full;
  wire                cpu_cmd_fire;
  wire                is_hit;
  reg                 is_hit_d1;
  wire                cpu_cmd_fire_1;
  wire                is_miss;
  wire                is_diff;
  reg                 flush_busy;
  reg                 flush_cnt_willIncrement;
  reg                 flush_cnt_willClear;
  reg        [3:0]    flush_cnt_valueNext;
  reg        [3:0]    flush_cnt_value;
  wire                flush_cnt_willOverflowIfInc;
  wire                flush_cnt_willOverflow;
  wire                flush_done;
  wire                cache_hit_gnt_0;
  wire                cache_hit_gnt_1;
  wire                cache_hit_gnt_2;
  wire                cache_hit_gnt_3;
  wire                cache_victim_gnt_0;
  wire                cache_victim_gnt_1;
  wire                cache_victim_gnt_2;
  wire                cache_victim_gnt_3;
  wire                cache_invld_gnt_0;
  wire                cache_invld_gnt_1;
  wire                cache_invld_gnt_2;
  wire                cache_invld_gnt_3;
  reg        [1:0]    evict_id_miss;
  wire       [53:0]   cpu_tag;
  wire       [3:0]    cpu_set;
  wire       [3:0]    cpu_bank_addr;
  wire       [3:0]    cpu_bank_index;
  wire                cpu_cmd_fire_2;
  reg        [63:0]   cpu_addr_d1;
  wire       [3:0]    cpu_set_d1;
  wire       [53:0]   cpu_tag_d1;
  wire       [3:0]    cpu_bank_addr_d1;
  wire       [3:0]    cpu_bank_index_d1;
  reg                 cpu_cmd_ready_1;
  wire       [511:0]  sram_banks_data_0;
  wire       [511:0]  sram_banks_data_1;
  wire       [511:0]  sram_banks_data_2;
  wire       [511:0]  sram_banks_data_3;
  wire                sram_banks_valid_0;
  wire                sram_banks_valid_1;
  wire                sram_banks_valid_2;
  wire                sram_banks_valid_3;
  reg                 next_level_cmd_valid_1;
  reg                 next_level_data_cnt_willIncrement;
  reg                 next_level_data_cnt_willClear;
  reg        [2:0]    next_level_data_cnt_valueNext;
  reg        [2:0]    next_level_data_cnt_value;
  wire                next_level_data_cnt_willOverflowIfInc;
  wire                next_level_data_cnt_willOverflow;
  wire       [3:0]    next_level_bank_addr;
  reg                 next_level_done;
  wire                when_ICache_l144;
  wire       [3:0]    _zz_cache_hit_gnt_0;
  wire       [3:0]    _zz_cache_hit_gnt_0_1;
  wire       [7:0]    _zz_cache_hit_gnt_0_2;
  wire       [7:0]    _zz_cache_hit_gnt_0_3;
  wire       [3:0]    _zz_cache_hit_gnt_0_4;
  wire       [3:0]    _zz_cache_invld_gnt_0;
  wire       [3:0]    _zz_cache_invld_gnt_0_1;
  wire       [7:0]    _zz_cache_invld_gnt_0_2;
  wire       [7:0]    _zz_cache_invld_gnt_0_3;
  wire       [3:0]    _zz_cache_invld_gnt_0_4;
  wire       [3:0]    _zz_cache_victim_gnt_0;
  wire       [3:0]    _zz_cache_victim_gnt_0_1;
  wire       [7:0]    _zz_cache_victim_gnt_0_2;
  wire       [7:0]    _zz_cache_victim_gnt_0_3;
  wire       [3:0]    _zz_cache_victim_gnt_0_4;
  wire                _zz_hit_id;
  wire                _zz_hit_id_1;
  wire                _zz_invld_id;
  wire                _zz_invld_id_1;
  wire                _zz_victim_id;
  wire                _zz_victim_id_1;
  wire       [15:0]   _zz_1;
  wire                _zz_2;
  wire                _zz_3;
  wire                _zz_4;
  wire                _zz_5;
  wire                _zz_6;
  wire                _zz_7;
  wire                _zz_8;
  wire                _zz_9;
  wire                _zz_10;
  wire                _zz_11;
  wire                _zz_12;
  wire                _zz_13;
  wire                _zz_14;
  wire                _zz_15;
  wire                _zz_16;
  wire                _zz_17;
  wire       [15:0]   _zz_18;
  wire                _zz_19;
  wire                _zz_20;
  wire                _zz_21;
  wire                _zz_22;
  wire                _zz_23;
  wire                _zz_24;
  wire                _zz_25;
  wire                _zz_26;
  wire                _zz_27;
  wire                _zz_28;
  wire                _zz_29;
  wire                _zz_30;
  wire                _zz_31;
  wire                _zz_32;
  wire                _zz_33;
  wire                _zz_34;
  wire                when_ICache_l176;
  reg        [15:0]   _zz_sram_0_ports_cmd_payload_wen;
  wire                when_ICache_l183;
  wire                when_ICache_l190;
  wire       [15:0]   _zz_35;
  wire                _zz_36;
  wire                _zz_37;
  wire                _zz_38;
  wire                _zz_39;
  wire                _zz_40;
  wire                _zz_41;
  wire                _zz_42;
  wire                _zz_43;
  wire                _zz_44;
  wire                _zz_45;
  wire                _zz_46;
  wire                _zz_47;
  wire                _zz_48;
  wire                _zz_49;
  wire                _zz_50;
  wire                _zz_51;
  wire                when_ICache_l212;
  wire                when_ICache_l219;
  wire                when_ICache_l222;
  wire                when_ICache_l227;
  wire                when_ICache_l232;
  wire                when_ICache_l235;
  wire       [15:0]   _zz_52;
  wire                _zz_53;
  wire                _zz_54;
  wire                _zz_55;
  wire                _zz_56;
  wire                _zz_57;
  wire                _zz_58;
  wire                _zz_59;
  wire                _zz_60;
  wire                _zz_61;
  wire                _zz_62;
  wire                _zz_63;
  wire                _zz_64;
  wire                _zz_65;
  wire                _zz_66;
  wire                _zz_67;
  wire                _zz_68;
  wire       [15:0]   _zz_69;
  wire                _zz_70;
  wire                _zz_71;
  wire                _zz_72;
  wire                _zz_73;
  wire                _zz_74;
  wire                _zz_75;
  wire                _zz_76;
  wire                _zz_77;
  wire                _zz_78;
  wire                _zz_79;
  wire                _zz_80;
  wire                _zz_81;
  wire                _zz_82;
  wire                _zz_83;
  wire                _zz_84;
  wire                _zz_85;
  wire                when_ICache_l176_1;
  reg        [15:0]   _zz_sram_1_ports_cmd_payload_wen;
  wire                when_ICache_l183_1;
  wire                when_ICache_l190_1;
  wire       [15:0]   _zz_86;
  wire                _zz_87;
  wire                _zz_88;
  wire                _zz_89;
  wire                _zz_90;
  wire                _zz_91;
  wire                _zz_92;
  wire                _zz_93;
  wire                _zz_94;
  wire                _zz_95;
  wire                _zz_96;
  wire                _zz_97;
  wire                _zz_98;
  wire                _zz_99;
  wire                _zz_100;
  wire                _zz_101;
  wire                _zz_102;
  wire                when_ICache_l212_1;
  wire                when_ICache_l219_1;
  wire                when_ICache_l222_1;
  wire                when_ICache_l227_1;
  wire                when_ICache_l232_1;
  wire                when_ICache_l235_1;
  wire       [15:0]   _zz_103;
  wire                _zz_104;
  wire                _zz_105;
  wire                _zz_106;
  wire                _zz_107;
  wire                _zz_108;
  wire                _zz_109;
  wire                _zz_110;
  wire                _zz_111;
  wire                _zz_112;
  wire                _zz_113;
  wire                _zz_114;
  wire                _zz_115;
  wire                _zz_116;
  wire                _zz_117;
  wire                _zz_118;
  wire                _zz_119;
  wire       [15:0]   _zz_120;
  wire                _zz_121;
  wire                _zz_122;
  wire                _zz_123;
  wire                _zz_124;
  wire                _zz_125;
  wire                _zz_126;
  wire                _zz_127;
  wire                _zz_128;
  wire                _zz_129;
  wire                _zz_130;
  wire                _zz_131;
  wire                _zz_132;
  wire                _zz_133;
  wire                _zz_134;
  wire                _zz_135;
  wire                _zz_136;
  wire                when_ICache_l176_2;
  reg        [15:0]   _zz_sram_2_ports_cmd_payload_wen;
  wire                when_ICache_l183_2;
  wire                when_ICache_l190_2;
  wire       [15:0]   _zz_137;
  wire                _zz_138;
  wire                _zz_139;
  wire                _zz_140;
  wire                _zz_141;
  wire                _zz_142;
  wire                _zz_143;
  wire                _zz_144;
  wire                _zz_145;
  wire                _zz_146;
  wire                _zz_147;
  wire                _zz_148;
  wire                _zz_149;
  wire                _zz_150;
  wire                _zz_151;
  wire                _zz_152;
  wire                _zz_153;
  wire                when_ICache_l212_2;
  wire                when_ICache_l219_2;
  wire                when_ICache_l222_2;
  wire                when_ICache_l227_2;
  wire                when_ICache_l232_2;
  wire                when_ICache_l235_2;
  wire       [15:0]   _zz_154;
  wire                _zz_155;
  wire                _zz_156;
  wire                _zz_157;
  wire                _zz_158;
  wire                _zz_159;
  wire                _zz_160;
  wire                _zz_161;
  wire                _zz_162;
  wire                _zz_163;
  wire                _zz_164;
  wire                _zz_165;
  wire                _zz_166;
  wire                _zz_167;
  wire                _zz_168;
  wire                _zz_169;
  wire                _zz_170;
  wire       [15:0]   _zz_171;
  wire                _zz_172;
  wire                _zz_173;
  wire                _zz_174;
  wire                _zz_175;
  wire                _zz_176;
  wire                _zz_177;
  wire                _zz_178;
  wire                _zz_179;
  wire                _zz_180;
  wire                _zz_181;
  wire                _zz_182;
  wire                _zz_183;
  wire                _zz_184;
  wire                _zz_185;
  wire                _zz_186;
  wire                _zz_187;
  wire                when_ICache_l176_3;
  reg        [15:0]   _zz_sram_3_ports_cmd_payload_wen;
  wire                when_ICache_l183_3;
  wire                when_ICache_l190_3;
  wire       [15:0]   _zz_188;
  wire                _zz_189;
  wire                _zz_190;
  wire                _zz_191;
  wire                _zz_192;
  wire                _zz_193;
  wire                _zz_194;
  wire                _zz_195;
  wire                _zz_196;
  wire                _zz_197;
  wire                _zz_198;
  wire                _zz_199;
  wire                _zz_200;
  wire                _zz_201;
  wire                _zz_202;
  wire                _zz_203;
  wire                _zz_204;
  wire                when_ICache_l212_3;
  wire                when_ICache_l219_3;
  wire                when_ICache_l222_3;
  wire                when_ICache_l227_3;
  wire                when_ICache_l232_3;
  wire                when_ICache_l235_3;
  wire       [511:0]  _zz_hit_data;
  wire       [31:0]   hit_data;
  wire       [511:0]  _zz_miss_data;
  wire       [31:0]   miss_data;
  function [15:0] zz__zz_sram_0_ports_cmd_payload_wen(input dummy);
    begin
      zz__zz_sram_0_ports_cmd_payload_wen = 16'h0;
      zz__zz_sram_0_ports_cmd_payload_wen[1] = 1'b1;
      zz__zz_sram_0_ports_cmd_payload_wen[0] = 1'b1;
    end
  endfunction
  wire [15:0] _zz_205;
  function [15:0] zz__zz_sram_1_ports_cmd_payload_wen(input dummy);
    begin
      zz__zz_sram_1_ports_cmd_payload_wen = 16'h0;
      zz__zz_sram_1_ports_cmd_payload_wen[1] = 1'b1;
      zz__zz_sram_1_ports_cmd_payload_wen[0] = 1'b1;
    end
  endfunction
  wire [15:0] _zz_206;
  function [15:0] zz__zz_sram_2_ports_cmd_payload_wen(input dummy);
    begin
      zz__zz_sram_2_ports_cmd_payload_wen = 16'h0;
      zz__zz_sram_2_ports_cmd_payload_wen[1] = 1'b1;
      zz__zz_sram_2_ports_cmd_payload_wen[0] = 1'b1;
    end
  endfunction
  wire [15:0] _zz_207;
  function [15:0] zz__zz_sram_3_ports_cmd_payload_wen(input dummy);
    begin
      zz__zz_sram_3_ports_cmd_payload_wen = 16'h0;
      zz__zz_sram_3_ports_cmd_payload_wen[1] = 1'b1;
      zz__zz_sram_3_ports_cmd_payload_wen[0] = 1'b1;
    end
  endfunction
  wire [15:0] _zz_208;

  assign _zz_flush_cnt_valueNext_1 = flush_cnt_willIncrement;
  assign _zz_flush_cnt_valueNext = {3'd0, _zz_flush_cnt_valueNext_1};
  assign _zz_next_level_data_cnt_valueNext_1 = next_level_data_cnt_willIncrement;
  assign _zz_next_level_data_cnt_valueNext = {2'd0, _zz_next_level_data_cnt_valueNext_1};
  assign _zz__zz_cache_hit_gnt_0_3 = (_zz_cache_hit_gnt_0_2 - _zz__zz_cache_hit_gnt_0_3_1);
  assign _zz__zz_cache_hit_gnt_0_3_2 = {_zz_cache_hit_gnt_0[3],{_zz_cache_hit_gnt_0[2],{_zz_cache_hit_gnt_0[1],_zz_cache_hit_gnt_0[0]}}};
  assign _zz__zz_cache_hit_gnt_0_3_1 = {4'd0, _zz__zz_cache_hit_gnt_0_3_2};
  assign _zz__zz_cache_invld_gnt_0_3 = (_zz_cache_invld_gnt_0_2 - _zz__zz_cache_invld_gnt_0_3_1);
  assign _zz__zz_cache_invld_gnt_0_3_2 = {_zz_cache_invld_gnt_0[3],{_zz_cache_invld_gnt_0[2],{_zz_cache_invld_gnt_0[1],_zz_cache_invld_gnt_0[0]}}};
  assign _zz__zz_cache_invld_gnt_0_3_1 = {4'd0, _zz__zz_cache_invld_gnt_0_3_2};
  assign _zz__zz_cache_victim_gnt_0_3 = (_zz_cache_victim_gnt_0_2 - _zz__zz_cache_victim_gnt_0_3_1);
  assign _zz__zz_cache_victim_gnt_0_3_2 = {_zz_cache_victim_gnt_0[3],{_zz_cache_victim_gnt_0[2],{_zz_cache_victim_gnt_0[1],_zz_cache_victim_gnt_0[0]}}};
  assign _zz__zz_cache_victim_gnt_0_3_1 = {4'd0, _zz__zz_cache_victim_gnt_0_3_2};
  assign _zz_sram_0_ports_cmd_payload_wen_1 = (next_level_data_cnt_value * 2'b10);
  assign _zz_sram_0_ports_cmd_payload_wdata = (next_level_data_cnt_value * 7'h40);
  assign _zz_sram_0_ports_cmd_payload_wstrb = (_zz_sram_0_ports_cmd_payload_wstrb_1 / 4'b1000);
  assign _zz_sram_0_ports_cmd_payload_wstrb_1 = (next_level_data_cnt_value * 7'h40);
  assign _zz_sram_1_ports_cmd_payload_wen_1 = (next_level_data_cnt_value * 2'b10);
  assign _zz_sram_1_ports_cmd_payload_wdata = (next_level_data_cnt_value * 7'h40);
  assign _zz_sram_1_ports_cmd_payload_wstrb = (_zz_sram_1_ports_cmd_payload_wstrb_1 / 4'b1000);
  assign _zz_sram_1_ports_cmd_payload_wstrb_1 = (next_level_data_cnt_value * 7'h40);
  assign _zz_sram_2_ports_cmd_payload_wen_1 = (next_level_data_cnt_value * 2'b10);
  assign _zz_sram_2_ports_cmd_payload_wdata = (next_level_data_cnt_value * 7'h40);
  assign _zz_sram_2_ports_cmd_payload_wstrb = (_zz_sram_2_ports_cmd_payload_wstrb_1 / 4'b1000);
  assign _zz_sram_2_ports_cmd_payload_wstrb_1 = (next_level_data_cnt_value * 7'h40);
  assign _zz_sram_3_ports_cmd_payload_wen_1 = (next_level_data_cnt_value * 2'b10);
  assign _zz_sram_3_ports_cmd_payload_wdata = (next_level_data_cnt_value * 7'h40);
  assign _zz_sram_3_ports_cmd_payload_wstrb = (_zz_sram_3_ports_cmd_payload_wstrb_1 / 4'b1000);
  assign _zz_sram_3_ports_cmd_payload_wstrb_1 = (next_level_data_cnt_value * 7'h40);
  always @(*) begin
    case(cpu_set)
      4'b0000 : begin
        _zz_cache_tag_0 = ways_0_metas_0_tag;
        _zz_cache_hit_0 = ways_0_metas_0_vld;
        _zz_cache_mru_0 = ways_0_metas_0_mru;
        _zz_cache_tag_1 = ways_1_metas_0_tag;
        _zz_cache_hit_1 = ways_1_metas_0_vld;
        _zz_cache_mru_1 = ways_1_metas_0_mru;
        _zz_cache_tag_2 = ways_2_metas_0_tag;
        _zz_cache_hit_2 = ways_2_metas_0_vld;
        _zz_cache_mru_2 = ways_2_metas_0_mru;
        _zz_cache_tag_3 = ways_3_metas_0_tag;
        _zz_cache_hit_3 = ways_3_metas_0_vld;
        _zz_cache_mru_3 = ways_3_metas_0_mru;
      end
      4'b0001 : begin
        _zz_cache_tag_0 = ways_0_metas_1_tag;
        _zz_cache_hit_0 = ways_0_metas_1_vld;
        _zz_cache_mru_0 = ways_0_metas_1_mru;
        _zz_cache_tag_1 = ways_1_metas_1_tag;
        _zz_cache_hit_1 = ways_1_metas_1_vld;
        _zz_cache_mru_1 = ways_1_metas_1_mru;
        _zz_cache_tag_2 = ways_2_metas_1_tag;
        _zz_cache_hit_2 = ways_2_metas_1_vld;
        _zz_cache_mru_2 = ways_2_metas_1_mru;
        _zz_cache_tag_3 = ways_3_metas_1_tag;
        _zz_cache_hit_3 = ways_3_metas_1_vld;
        _zz_cache_mru_3 = ways_3_metas_1_mru;
      end
      4'b0010 : begin
        _zz_cache_tag_0 = ways_0_metas_2_tag;
        _zz_cache_hit_0 = ways_0_metas_2_vld;
        _zz_cache_mru_0 = ways_0_metas_2_mru;
        _zz_cache_tag_1 = ways_1_metas_2_tag;
        _zz_cache_hit_1 = ways_1_metas_2_vld;
        _zz_cache_mru_1 = ways_1_metas_2_mru;
        _zz_cache_tag_2 = ways_2_metas_2_tag;
        _zz_cache_hit_2 = ways_2_metas_2_vld;
        _zz_cache_mru_2 = ways_2_metas_2_mru;
        _zz_cache_tag_3 = ways_3_metas_2_tag;
        _zz_cache_hit_3 = ways_3_metas_2_vld;
        _zz_cache_mru_3 = ways_3_metas_2_mru;
      end
      4'b0011 : begin
        _zz_cache_tag_0 = ways_0_metas_3_tag;
        _zz_cache_hit_0 = ways_0_metas_3_vld;
        _zz_cache_mru_0 = ways_0_metas_3_mru;
        _zz_cache_tag_1 = ways_1_metas_3_tag;
        _zz_cache_hit_1 = ways_1_metas_3_vld;
        _zz_cache_mru_1 = ways_1_metas_3_mru;
        _zz_cache_tag_2 = ways_2_metas_3_tag;
        _zz_cache_hit_2 = ways_2_metas_3_vld;
        _zz_cache_mru_2 = ways_2_metas_3_mru;
        _zz_cache_tag_3 = ways_3_metas_3_tag;
        _zz_cache_hit_3 = ways_3_metas_3_vld;
        _zz_cache_mru_3 = ways_3_metas_3_mru;
      end
      4'b0100 : begin
        _zz_cache_tag_0 = ways_0_metas_4_tag;
        _zz_cache_hit_0 = ways_0_metas_4_vld;
        _zz_cache_mru_0 = ways_0_metas_4_mru;
        _zz_cache_tag_1 = ways_1_metas_4_tag;
        _zz_cache_hit_1 = ways_1_metas_4_vld;
        _zz_cache_mru_1 = ways_1_metas_4_mru;
        _zz_cache_tag_2 = ways_2_metas_4_tag;
        _zz_cache_hit_2 = ways_2_metas_4_vld;
        _zz_cache_mru_2 = ways_2_metas_4_mru;
        _zz_cache_tag_3 = ways_3_metas_4_tag;
        _zz_cache_hit_3 = ways_3_metas_4_vld;
        _zz_cache_mru_3 = ways_3_metas_4_mru;
      end
      4'b0101 : begin
        _zz_cache_tag_0 = ways_0_metas_5_tag;
        _zz_cache_hit_0 = ways_0_metas_5_vld;
        _zz_cache_mru_0 = ways_0_metas_5_mru;
        _zz_cache_tag_1 = ways_1_metas_5_tag;
        _zz_cache_hit_1 = ways_1_metas_5_vld;
        _zz_cache_mru_1 = ways_1_metas_5_mru;
        _zz_cache_tag_2 = ways_2_metas_5_tag;
        _zz_cache_hit_2 = ways_2_metas_5_vld;
        _zz_cache_mru_2 = ways_2_metas_5_mru;
        _zz_cache_tag_3 = ways_3_metas_5_tag;
        _zz_cache_hit_3 = ways_3_metas_5_vld;
        _zz_cache_mru_3 = ways_3_metas_5_mru;
      end
      4'b0110 : begin
        _zz_cache_tag_0 = ways_0_metas_6_tag;
        _zz_cache_hit_0 = ways_0_metas_6_vld;
        _zz_cache_mru_0 = ways_0_metas_6_mru;
        _zz_cache_tag_1 = ways_1_metas_6_tag;
        _zz_cache_hit_1 = ways_1_metas_6_vld;
        _zz_cache_mru_1 = ways_1_metas_6_mru;
        _zz_cache_tag_2 = ways_2_metas_6_tag;
        _zz_cache_hit_2 = ways_2_metas_6_vld;
        _zz_cache_mru_2 = ways_2_metas_6_mru;
        _zz_cache_tag_3 = ways_3_metas_6_tag;
        _zz_cache_hit_3 = ways_3_metas_6_vld;
        _zz_cache_mru_3 = ways_3_metas_6_mru;
      end
      4'b0111 : begin
        _zz_cache_tag_0 = ways_0_metas_7_tag;
        _zz_cache_hit_0 = ways_0_metas_7_vld;
        _zz_cache_mru_0 = ways_0_metas_7_mru;
        _zz_cache_tag_1 = ways_1_metas_7_tag;
        _zz_cache_hit_1 = ways_1_metas_7_vld;
        _zz_cache_mru_1 = ways_1_metas_7_mru;
        _zz_cache_tag_2 = ways_2_metas_7_tag;
        _zz_cache_hit_2 = ways_2_metas_7_vld;
        _zz_cache_mru_2 = ways_2_metas_7_mru;
        _zz_cache_tag_3 = ways_3_metas_7_tag;
        _zz_cache_hit_3 = ways_3_metas_7_vld;
        _zz_cache_mru_3 = ways_3_metas_7_mru;
      end
      4'b1000 : begin
        _zz_cache_tag_0 = ways_0_metas_8_tag;
        _zz_cache_hit_0 = ways_0_metas_8_vld;
        _zz_cache_mru_0 = ways_0_metas_8_mru;
        _zz_cache_tag_1 = ways_1_metas_8_tag;
        _zz_cache_hit_1 = ways_1_metas_8_vld;
        _zz_cache_mru_1 = ways_1_metas_8_mru;
        _zz_cache_tag_2 = ways_2_metas_8_tag;
        _zz_cache_hit_2 = ways_2_metas_8_vld;
        _zz_cache_mru_2 = ways_2_metas_8_mru;
        _zz_cache_tag_3 = ways_3_metas_8_tag;
        _zz_cache_hit_3 = ways_3_metas_8_vld;
        _zz_cache_mru_3 = ways_3_metas_8_mru;
      end
      4'b1001 : begin
        _zz_cache_tag_0 = ways_0_metas_9_tag;
        _zz_cache_hit_0 = ways_0_metas_9_vld;
        _zz_cache_mru_0 = ways_0_metas_9_mru;
        _zz_cache_tag_1 = ways_1_metas_9_tag;
        _zz_cache_hit_1 = ways_1_metas_9_vld;
        _zz_cache_mru_1 = ways_1_metas_9_mru;
        _zz_cache_tag_2 = ways_2_metas_9_tag;
        _zz_cache_hit_2 = ways_2_metas_9_vld;
        _zz_cache_mru_2 = ways_2_metas_9_mru;
        _zz_cache_tag_3 = ways_3_metas_9_tag;
        _zz_cache_hit_3 = ways_3_metas_9_vld;
        _zz_cache_mru_3 = ways_3_metas_9_mru;
      end
      4'b1010 : begin
        _zz_cache_tag_0 = ways_0_metas_10_tag;
        _zz_cache_hit_0 = ways_0_metas_10_vld;
        _zz_cache_mru_0 = ways_0_metas_10_mru;
        _zz_cache_tag_1 = ways_1_metas_10_tag;
        _zz_cache_hit_1 = ways_1_metas_10_vld;
        _zz_cache_mru_1 = ways_1_metas_10_mru;
        _zz_cache_tag_2 = ways_2_metas_10_tag;
        _zz_cache_hit_2 = ways_2_metas_10_vld;
        _zz_cache_mru_2 = ways_2_metas_10_mru;
        _zz_cache_tag_3 = ways_3_metas_10_tag;
        _zz_cache_hit_3 = ways_3_metas_10_vld;
        _zz_cache_mru_3 = ways_3_metas_10_mru;
      end
      4'b1011 : begin
        _zz_cache_tag_0 = ways_0_metas_11_tag;
        _zz_cache_hit_0 = ways_0_metas_11_vld;
        _zz_cache_mru_0 = ways_0_metas_11_mru;
        _zz_cache_tag_1 = ways_1_metas_11_tag;
        _zz_cache_hit_1 = ways_1_metas_11_vld;
        _zz_cache_mru_1 = ways_1_metas_11_mru;
        _zz_cache_tag_2 = ways_2_metas_11_tag;
        _zz_cache_hit_2 = ways_2_metas_11_vld;
        _zz_cache_mru_2 = ways_2_metas_11_mru;
        _zz_cache_tag_3 = ways_3_metas_11_tag;
        _zz_cache_hit_3 = ways_3_metas_11_vld;
        _zz_cache_mru_3 = ways_3_metas_11_mru;
      end
      4'b1100 : begin
        _zz_cache_tag_0 = ways_0_metas_12_tag;
        _zz_cache_hit_0 = ways_0_metas_12_vld;
        _zz_cache_mru_0 = ways_0_metas_12_mru;
        _zz_cache_tag_1 = ways_1_metas_12_tag;
        _zz_cache_hit_1 = ways_1_metas_12_vld;
        _zz_cache_mru_1 = ways_1_metas_12_mru;
        _zz_cache_tag_2 = ways_2_metas_12_tag;
        _zz_cache_hit_2 = ways_2_metas_12_vld;
        _zz_cache_mru_2 = ways_2_metas_12_mru;
        _zz_cache_tag_3 = ways_3_metas_12_tag;
        _zz_cache_hit_3 = ways_3_metas_12_vld;
        _zz_cache_mru_3 = ways_3_metas_12_mru;
      end
      4'b1101 : begin
        _zz_cache_tag_0 = ways_0_metas_13_tag;
        _zz_cache_hit_0 = ways_0_metas_13_vld;
        _zz_cache_mru_0 = ways_0_metas_13_mru;
        _zz_cache_tag_1 = ways_1_metas_13_tag;
        _zz_cache_hit_1 = ways_1_metas_13_vld;
        _zz_cache_mru_1 = ways_1_metas_13_mru;
        _zz_cache_tag_2 = ways_2_metas_13_tag;
        _zz_cache_hit_2 = ways_2_metas_13_vld;
        _zz_cache_mru_2 = ways_2_metas_13_mru;
        _zz_cache_tag_3 = ways_3_metas_13_tag;
        _zz_cache_hit_3 = ways_3_metas_13_vld;
        _zz_cache_mru_3 = ways_3_metas_13_mru;
      end
      4'b1110 : begin
        _zz_cache_tag_0 = ways_0_metas_14_tag;
        _zz_cache_hit_0 = ways_0_metas_14_vld;
        _zz_cache_mru_0 = ways_0_metas_14_mru;
        _zz_cache_tag_1 = ways_1_metas_14_tag;
        _zz_cache_hit_1 = ways_1_metas_14_vld;
        _zz_cache_mru_1 = ways_1_metas_14_mru;
        _zz_cache_tag_2 = ways_2_metas_14_tag;
        _zz_cache_hit_2 = ways_2_metas_14_vld;
        _zz_cache_mru_2 = ways_2_metas_14_mru;
        _zz_cache_tag_3 = ways_3_metas_14_tag;
        _zz_cache_hit_3 = ways_3_metas_14_vld;
        _zz_cache_mru_3 = ways_3_metas_14_mru;
      end
      default : begin
        _zz_cache_tag_0 = ways_0_metas_15_tag;
        _zz_cache_hit_0 = ways_0_metas_15_vld;
        _zz_cache_mru_0 = ways_0_metas_15_mru;
        _zz_cache_tag_1 = ways_1_metas_15_tag;
        _zz_cache_hit_1 = ways_1_metas_15_vld;
        _zz_cache_mru_1 = ways_1_metas_15_mru;
        _zz_cache_tag_2 = ways_2_metas_15_tag;
        _zz_cache_hit_2 = ways_2_metas_15_vld;
        _zz_cache_mru_2 = ways_2_metas_15_mru;
        _zz_cache_tag_3 = ways_3_metas_15_tag;
        _zz_cache_hit_3 = ways_3_metas_15_vld;
        _zz_cache_mru_3 = ways_3_metas_15_mru;
      end
    endcase
  end

  always @(*) begin
    case(cpu_set_d1)
      4'b0000 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_0_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_0_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_0_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_0_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_0_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_0_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_0_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_0_mru;
      end
      4'b0001 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_1_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_1_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_1_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_1_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_1_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_1_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_1_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_1_mru;
      end
      4'b0010 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_2_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_2_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_2_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_2_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_2_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_2_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_2_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_2_mru;
      end
      4'b0011 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_3_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_3_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_3_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_3_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_3_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_3_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_3_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_3_mru;
      end
      4'b0100 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_4_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_4_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_4_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_4_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_4_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_4_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_4_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_4_mru;
      end
      4'b0101 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_5_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_5_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_5_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_5_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_5_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_5_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_5_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_5_mru;
      end
      4'b0110 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_6_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_6_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_6_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_6_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_6_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_6_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_6_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_6_mru;
      end
      4'b0111 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_7_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_7_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_7_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_7_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_7_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_7_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_7_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_7_mru;
      end
      4'b1000 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_8_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_8_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_8_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_8_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_8_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_8_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_8_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_8_mru;
      end
      4'b1001 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_9_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_9_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_9_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_9_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_9_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_9_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_9_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_9_mru;
      end
      4'b1010 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_10_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_10_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_10_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_10_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_10_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_10_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_10_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_10_mru;
      end
      4'b1011 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_11_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_11_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_11_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_11_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_11_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_11_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_11_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_11_mru;
      end
      4'b1100 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_12_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_12_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_12_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_12_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_12_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_12_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_12_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_12_mru;
      end
      4'b1101 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_13_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_13_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_13_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_13_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_13_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_13_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_13_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_13_mru;
      end
      4'b1110 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_14_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_14_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_14_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_14_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_14_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_14_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_14_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_14_mru;
      end
      default : begin
        _zz_cache_invld_d1_0 = ways_0_metas_15_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_15_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_15_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_15_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_15_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_15_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_15_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_15_mru;
      end
    endcase
  end

  always @(*) begin
    case(hit_id_d1)
      2'b00 : begin
        _zz__zz_hit_data = sram_banks_data_0;
        _zz_cpu_rsp_valid = sram_banks_valid_0;
      end
      2'b01 : begin
        _zz__zz_hit_data = sram_banks_data_1;
        _zz_cpu_rsp_valid = sram_banks_valid_1;
      end
      2'b10 : begin
        _zz__zz_hit_data = sram_banks_data_2;
        _zz_cpu_rsp_valid = sram_banks_valid_2;
      end
      default : begin
        _zz__zz_hit_data = sram_banks_data_3;
        _zz_cpu_rsp_valid = sram_banks_valid_3;
      end
    endcase
  end

  always @(*) begin
    case(cpu_bank_index_d1)
      4'b0000 : begin
        _zz_hit_data_1 = _zz_hit_data[31 : 0];
        _zz_miss_data_1 = _zz_miss_data[31 : 0];
      end
      4'b0001 : begin
        _zz_hit_data_1 = _zz_hit_data[63 : 32];
        _zz_miss_data_1 = _zz_miss_data[63 : 32];
      end
      4'b0010 : begin
        _zz_hit_data_1 = _zz_hit_data[95 : 64];
        _zz_miss_data_1 = _zz_miss_data[95 : 64];
      end
      4'b0011 : begin
        _zz_hit_data_1 = _zz_hit_data[127 : 96];
        _zz_miss_data_1 = _zz_miss_data[127 : 96];
      end
      4'b0100 : begin
        _zz_hit_data_1 = _zz_hit_data[159 : 128];
        _zz_miss_data_1 = _zz_miss_data[159 : 128];
      end
      4'b0101 : begin
        _zz_hit_data_1 = _zz_hit_data[191 : 160];
        _zz_miss_data_1 = _zz_miss_data[191 : 160];
      end
      4'b0110 : begin
        _zz_hit_data_1 = _zz_hit_data[223 : 192];
        _zz_miss_data_1 = _zz_miss_data[223 : 192];
      end
      4'b0111 : begin
        _zz_hit_data_1 = _zz_hit_data[255 : 224];
        _zz_miss_data_1 = _zz_miss_data[255 : 224];
      end
      4'b1000 : begin
        _zz_hit_data_1 = _zz_hit_data[287 : 256];
        _zz_miss_data_1 = _zz_miss_data[287 : 256];
      end
      4'b1001 : begin
        _zz_hit_data_1 = _zz_hit_data[319 : 288];
        _zz_miss_data_1 = _zz_miss_data[319 : 288];
      end
      4'b1010 : begin
        _zz_hit_data_1 = _zz_hit_data[351 : 320];
        _zz_miss_data_1 = _zz_miss_data[351 : 320];
      end
      4'b1011 : begin
        _zz_hit_data_1 = _zz_hit_data[383 : 352];
        _zz_miss_data_1 = _zz_miss_data[383 : 352];
      end
      4'b1100 : begin
        _zz_hit_data_1 = _zz_hit_data[415 : 384];
        _zz_miss_data_1 = _zz_miss_data[415 : 384];
      end
      4'b1101 : begin
        _zz_hit_data_1 = _zz_hit_data[447 : 416];
        _zz_miss_data_1 = _zz_miss_data[447 : 416];
      end
      4'b1110 : begin
        _zz_hit_data_1 = _zz_hit_data[479 : 448];
        _zz_miss_data_1 = _zz_miss_data[479 : 448];
      end
      default : begin
        _zz_hit_data_1 = _zz_hit_data[511 : 480];
        _zz_miss_data_1 = _zz_miss_data[511 : 480];
      end
    endcase
  end

  always @(*) begin
    case(evict_id_miss)
      2'b00 : begin
        _zz__zz_miss_data = sram_banks_data_0;
        _zz_cpu_rsp_valid_1 = sram_banks_valid_0;
      end
      2'b01 : begin
        _zz__zz_miss_data = sram_banks_data_1;
        _zz_cpu_rsp_valid_1 = sram_banks_valid_1;
      end
      2'b10 : begin
        _zz__zz_miss_data = sram_banks_data_2;
        _zz_cpu_rsp_valid_1 = sram_banks_valid_2;
      end
      default : begin
        _zz__zz_miss_data = sram_banks_data_3;
        _zz_cpu_rsp_valid_1 = sram_banks_valid_3;
      end
    endcase
  end

  assign mru_full = (&{cache_mru_3,{cache_mru_2,{cache_mru_1,cache_mru_0}}});
  assign cpu_cmd_fire = (cpu_cmd_valid && cpu_cmd_ready);
  assign is_hit = ((|{cache_hit_3,{cache_hit_2,{cache_hit_1,cache_hit_0}}}) && cpu_cmd_fire);
  assign cpu_cmd_fire_1 = (cpu_cmd_valid && cpu_cmd_ready);
  assign is_miss = ((! (|{cache_hit_3,{cache_hit_2,{cache_hit_1,cache_hit_0}}})) && cpu_cmd_fire_1);
  assign is_diff = (! (|{cache_victim_3,{cache_victim_2,{cache_victim_1,cache_victim_0}}}));
  always @(*) begin
    flush_cnt_willIncrement = 1'b0;
    if(!when_ICache_l144) begin
      if(flush_busy) begin
        flush_cnt_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    flush_cnt_willClear = 1'b0;
    if(when_ICache_l144) begin
      flush_cnt_willClear = 1'b1;
    end
  end

  assign flush_cnt_willOverflowIfInc = (flush_cnt_value == 4'b1111);
  assign flush_cnt_willOverflow = (flush_cnt_willOverflowIfInc && flush_cnt_willIncrement);
  always @(*) begin
    flush_cnt_valueNext = (flush_cnt_value + _zz_flush_cnt_valueNext);
    if(flush_cnt_willClear) begin
      flush_cnt_valueNext = 4'b0000;
    end
  end

  assign flush_done = (flush_busy && (flush_cnt_value == 4'b1111));
  assign cpu_tag = cpu_cmd_payload_addr[63 : 10];
  assign cpu_set = cpu_cmd_payload_addr[9 : 6];
  assign cpu_bank_addr = cpu_cmd_payload_addr[9 : 6];
  assign cpu_bank_index = cpu_cmd_payload_addr[5 : 2];
  assign cpu_cmd_fire_2 = (cpu_cmd_valid && cpu_cmd_ready);
  assign cpu_set_d1 = cpu_addr_d1[9 : 6];
  assign cpu_tag_d1 = cpu_addr_d1[63 : 10];
  assign cpu_bank_addr_d1 = cpu_addr_d1[9 : 6];
  assign cpu_bank_index_d1 = cpu_addr_d1[5 : 2];
  always @(*) begin
    next_level_data_cnt_willIncrement = 1'b0;
    if(!is_miss) begin
      if(!next_level_done) begin
        if(next_level_rsp_valid) begin
          next_level_data_cnt_willIncrement = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    next_level_data_cnt_willClear = 1'b0;
    if(is_miss) begin
      next_level_data_cnt_willClear = 1'b1;
    end else begin
      if(next_level_done) begin
        next_level_data_cnt_willClear = 1'b1;
      end
    end
  end

  assign next_level_data_cnt_willOverflowIfInc = (next_level_data_cnt_value == 3'b111);
  assign next_level_data_cnt_willOverflow = (next_level_data_cnt_willOverflowIfInc && next_level_data_cnt_willIncrement);
  always @(*) begin
    next_level_data_cnt_valueNext = (next_level_data_cnt_value + _zz_next_level_data_cnt_valueNext);
    if(next_level_data_cnt_willClear) begin
      next_level_data_cnt_valueNext = 3'b000;
    end
  end

  assign next_level_bank_addr = cpu_addr_d1[9 : 6];
  assign when_ICache_l144 = (flush_busy && (flush_cnt_value == 4'b1111));
  assign _zz_cache_hit_gnt_0 = 4'b0001;
  assign _zz_cache_hit_gnt_0_1 = {cache_hit_3,{cache_hit_2,{cache_hit_1,cache_hit_0}}};
  assign _zz_cache_hit_gnt_0_2 = {_zz_cache_hit_gnt_0_1,_zz_cache_hit_gnt_0_1};
  assign _zz_cache_hit_gnt_0_3 = (_zz_cache_hit_gnt_0_2 & (~ _zz__zz_cache_hit_gnt_0_3));
  assign _zz_cache_hit_gnt_0_4 = (_zz_cache_hit_gnt_0_3[7 : 4] | _zz_cache_hit_gnt_0_3[3 : 0]);
  assign cache_hit_gnt_0 = _zz_cache_hit_gnt_0_4[0];
  assign cache_hit_gnt_1 = _zz_cache_hit_gnt_0_4[1];
  assign cache_hit_gnt_2 = _zz_cache_hit_gnt_0_4[2];
  assign cache_hit_gnt_3 = _zz_cache_hit_gnt_0_4[3];
  assign _zz_cache_invld_gnt_0 = 4'b0001;
  assign _zz_cache_invld_gnt_0_1 = {cache_invld_d1_3,{cache_invld_d1_2,{cache_invld_d1_1,cache_invld_d1_0}}};
  assign _zz_cache_invld_gnt_0_2 = {_zz_cache_invld_gnt_0_1,_zz_cache_invld_gnt_0_1};
  assign _zz_cache_invld_gnt_0_3 = (_zz_cache_invld_gnt_0_2 & (~ _zz__zz_cache_invld_gnt_0_3));
  assign _zz_cache_invld_gnt_0_4 = (_zz_cache_invld_gnt_0_3[7 : 4] | _zz_cache_invld_gnt_0_3[3 : 0]);
  assign cache_invld_gnt_0 = _zz_cache_invld_gnt_0_4[0];
  assign cache_invld_gnt_1 = _zz_cache_invld_gnt_0_4[1];
  assign cache_invld_gnt_2 = _zz_cache_invld_gnt_0_4[2];
  assign cache_invld_gnt_3 = _zz_cache_invld_gnt_0_4[3];
  assign _zz_cache_victim_gnt_0 = 4'b0001;
  assign _zz_cache_victim_gnt_0_1 = {cache_victim_3,{cache_victim_2,{cache_victim_1,cache_victim_0}}};
  assign _zz_cache_victim_gnt_0_2 = {_zz_cache_victim_gnt_0_1,_zz_cache_victim_gnt_0_1};
  assign _zz_cache_victim_gnt_0_3 = (_zz_cache_victim_gnt_0_2 & (~ _zz__zz_cache_victim_gnt_0_3));
  assign _zz_cache_victim_gnt_0_4 = (_zz_cache_victim_gnt_0_3[7 : 4] | _zz_cache_victim_gnt_0_3[3 : 0]);
  assign cache_victim_gnt_0 = _zz_cache_victim_gnt_0_4[0];
  assign cache_victim_gnt_1 = _zz_cache_victim_gnt_0_4[1];
  assign cache_victim_gnt_2 = _zz_cache_victim_gnt_0_4[2];
  assign cache_victim_gnt_3 = _zz_cache_victim_gnt_0_4[3];
  assign _zz_hit_id = (cache_hit_gnt_1 || cache_hit_gnt_3);
  assign _zz_hit_id_1 = (cache_hit_gnt_2 || cache_hit_gnt_3);
  assign hit_id = {_zz_hit_id_1,_zz_hit_id};
  assign _zz_invld_id = (cache_invld_gnt_1 || cache_invld_gnt_3);
  assign _zz_invld_id_1 = (cache_invld_gnt_2 || cache_invld_gnt_3);
  assign invld_id = {_zz_invld_id_1,_zz_invld_id};
  assign _zz_victim_id = (cache_victim_gnt_1 || cache_victim_gnt_3);
  assign _zz_victim_id_1 = (cache_victim_gnt_2 || cache_victim_gnt_3);
  assign victim_id = {_zz_victim_id_1,_zz_victim_id};
  assign evict_id = (is_diff ? invld_id : victim_id);
  assign _zz_1 = ({15'd0,1'b1} <<< cpu_set);
  assign _zz_2 = _zz_1[0];
  assign _zz_3 = _zz_1[1];
  assign _zz_4 = _zz_1[2];
  assign _zz_5 = _zz_1[3];
  assign _zz_6 = _zz_1[4];
  assign _zz_7 = _zz_1[5];
  assign _zz_8 = _zz_1[6];
  assign _zz_9 = _zz_1[7];
  assign _zz_10 = _zz_1[8];
  assign _zz_11 = _zz_1[9];
  assign _zz_12 = _zz_1[10];
  assign _zz_13 = _zz_1[11];
  assign _zz_14 = _zz_1[12];
  assign _zz_15 = _zz_1[13];
  assign _zz_16 = _zz_1[14];
  assign _zz_17 = _zz_1[15];
  assign cache_tag_0 = _zz_cache_tag_0;
  assign cache_hit_0 = ((cache_tag_0 == cpu_tag) && _zz_cache_hit_0);
  assign cache_mru_0 = _zz_cache_mru_0;
  assign _zz_18 = ({15'd0,1'b1} <<< cpu_set_d1);
  assign _zz_19 = _zz_18[0];
  assign _zz_20 = _zz_18[1];
  assign _zz_21 = _zz_18[2];
  assign _zz_22 = _zz_18[3];
  assign _zz_23 = _zz_18[4];
  assign _zz_24 = _zz_18[5];
  assign _zz_25 = _zz_18[6];
  assign _zz_26 = _zz_18[7];
  assign _zz_27 = _zz_18[8];
  assign _zz_28 = _zz_18[9];
  assign _zz_29 = _zz_18[10];
  assign _zz_30 = _zz_18[11];
  assign _zz_31 = _zz_18[12];
  assign _zz_32 = _zz_18[13];
  assign _zz_33 = _zz_18[14];
  assign _zz_34 = _zz_18[15];
  assign cache_invld_d1_0 = (! _zz_cache_invld_d1_0);
  assign cache_lru_d1_0 = (! _zz_cache_lru_d1_0);
  assign cache_victim_0 = (cache_invld_d1_0 && cache_lru_d1_0);
  assign sram_banks_data_0 = sram_0_ports_rsp_payload_data;
  assign sram_banks_valid_0 = sram_0_ports_rsp_valid;
  assign when_ICache_l176 = (is_hit && (2'b00 == hit_id));
  always @(*) begin
    if(when_ICache_l176) begin
      sram_0_ports_cmd_payload_addr = cpu_bank_addr;
    end else begin
      if(when_ICache_l183) begin
        sram_0_ports_cmd_payload_addr = cpu_bank_addr_d1;
      end else begin
        if(when_ICache_l190) begin
          sram_0_ports_cmd_payload_addr = next_level_bank_addr;
        end else begin
          sram_0_ports_cmd_payload_addr = 4'b0000;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l176) begin
      sram_0_ports_cmd_valid = 1'b1;
    end else begin
      if(when_ICache_l183) begin
        sram_0_ports_cmd_valid = 1'b1;
      end else begin
        if(when_ICache_l190) begin
          sram_0_ports_cmd_valid = 1'b1;
        end else begin
          sram_0_ports_cmd_valid = 1'b0;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l176) begin
      sram_0_ports_cmd_payload_wen = 16'h0;
    end else begin
      if(when_ICache_l183) begin
        sram_0_ports_cmd_payload_wen = 16'h0;
      end else begin
        if(when_ICache_l190) begin
          sram_0_ports_cmd_payload_wen = (_zz_sram_0_ports_cmd_payload_wen <<< _zz_sram_0_ports_cmd_payload_wen_1);
        end else begin
          sram_0_ports_cmd_payload_wen = 16'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l176) begin
      sram_0_ports_cmd_payload_wdata = 512'h0;
    end else begin
      if(when_ICache_l183) begin
        sram_0_ports_cmd_payload_wdata = 512'h0;
      end else begin
        if(when_ICache_l190) begin
          sram_0_ports_cmd_payload_wdata = ({448'h0,next_level_rsp_payload_data} <<< _zz_sram_0_ports_cmd_payload_wdata);
        end else begin
          sram_0_ports_cmd_payload_wdata = 512'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l176) begin
      sram_0_ports_cmd_payload_wstrb = 64'h0;
    end else begin
      if(when_ICache_l183) begin
        sram_0_ports_cmd_payload_wstrb = 64'h0;
      end else begin
        if(when_ICache_l190) begin
          sram_0_ports_cmd_payload_wstrb = ({56'h0,8'hff} <<< _zz_sram_0_ports_cmd_payload_wstrb);
        end else begin
          sram_0_ports_cmd_payload_wstrb = 64'h0;
        end
      end
    end
  end

  assign _zz_205 = zz__zz_sram_0_ports_cmd_payload_wen(1'b0);
  always @(*) _zz_sram_0_ports_cmd_payload_wen = _zz_205;
  assign when_ICache_l183 = (next_level_done && (2'b00 == evict_id_miss));
  assign when_ICache_l190 = (next_level_rsp_valid && (2'b00 == evict_id_miss));
  assign _zz_35 = ({15'd0,1'b1} <<< flush_cnt_value);
  assign _zz_36 = _zz_35[0];
  assign _zz_37 = _zz_35[1];
  assign _zz_38 = _zz_35[2];
  assign _zz_39 = _zz_35[3];
  assign _zz_40 = _zz_35[4];
  assign _zz_41 = _zz_35[5];
  assign _zz_42 = _zz_35[6];
  assign _zz_43 = _zz_35[7];
  assign _zz_44 = _zz_35[8];
  assign _zz_45 = _zz_35[9];
  assign _zz_46 = _zz_35[10];
  assign _zz_47 = _zz_35[11];
  assign _zz_48 = _zz_35[12];
  assign _zz_49 = _zz_35[13];
  assign _zz_50 = _zz_35[14];
  assign _zz_51 = _zz_35[15];
  assign when_ICache_l212 = (is_hit && mru_full);
  assign when_ICache_l219 = (is_hit && cache_hit_0);
  assign when_ICache_l222 = (next_level_done && (2'b00 == evict_id_miss));
  assign when_ICache_l227 = (next_level_done && (2'b00 == evict_id_miss));
  assign when_ICache_l232 = (flush || is_miss);
  assign when_ICache_l235 = (flush_done || next_level_done);
  assign _zz_52 = ({15'd0,1'b1} <<< cpu_set);
  assign _zz_53 = _zz_52[0];
  assign _zz_54 = _zz_52[1];
  assign _zz_55 = _zz_52[2];
  assign _zz_56 = _zz_52[3];
  assign _zz_57 = _zz_52[4];
  assign _zz_58 = _zz_52[5];
  assign _zz_59 = _zz_52[6];
  assign _zz_60 = _zz_52[7];
  assign _zz_61 = _zz_52[8];
  assign _zz_62 = _zz_52[9];
  assign _zz_63 = _zz_52[10];
  assign _zz_64 = _zz_52[11];
  assign _zz_65 = _zz_52[12];
  assign _zz_66 = _zz_52[13];
  assign _zz_67 = _zz_52[14];
  assign _zz_68 = _zz_52[15];
  assign cache_tag_1 = _zz_cache_tag_1;
  assign cache_hit_1 = ((cache_tag_1 == cpu_tag) && _zz_cache_hit_1);
  assign cache_mru_1 = _zz_cache_mru_1;
  assign _zz_69 = ({15'd0,1'b1} <<< cpu_set_d1);
  assign _zz_70 = _zz_69[0];
  assign _zz_71 = _zz_69[1];
  assign _zz_72 = _zz_69[2];
  assign _zz_73 = _zz_69[3];
  assign _zz_74 = _zz_69[4];
  assign _zz_75 = _zz_69[5];
  assign _zz_76 = _zz_69[6];
  assign _zz_77 = _zz_69[7];
  assign _zz_78 = _zz_69[8];
  assign _zz_79 = _zz_69[9];
  assign _zz_80 = _zz_69[10];
  assign _zz_81 = _zz_69[11];
  assign _zz_82 = _zz_69[12];
  assign _zz_83 = _zz_69[13];
  assign _zz_84 = _zz_69[14];
  assign _zz_85 = _zz_69[15];
  assign cache_invld_d1_1 = (! _zz_cache_invld_d1_1);
  assign cache_lru_d1_1 = (! _zz_cache_lru_d1_1);
  assign cache_victim_1 = (cache_invld_d1_1 && cache_lru_d1_1);
  assign sram_banks_data_1 = sram_1_ports_rsp_payload_data;
  assign sram_banks_valid_1 = sram_1_ports_rsp_valid;
  assign when_ICache_l176_1 = (is_hit && (2'b01 == hit_id));
  always @(*) begin
    if(when_ICache_l176_1) begin
      sram_1_ports_cmd_payload_addr = cpu_bank_addr;
    end else begin
      if(when_ICache_l183_1) begin
        sram_1_ports_cmd_payload_addr = cpu_bank_addr_d1;
      end else begin
        if(when_ICache_l190_1) begin
          sram_1_ports_cmd_payload_addr = next_level_bank_addr;
        end else begin
          sram_1_ports_cmd_payload_addr = 4'b0000;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l176_1) begin
      sram_1_ports_cmd_valid = 1'b1;
    end else begin
      if(when_ICache_l183_1) begin
        sram_1_ports_cmd_valid = 1'b1;
      end else begin
        if(when_ICache_l190_1) begin
          sram_1_ports_cmd_valid = 1'b1;
        end else begin
          sram_1_ports_cmd_valid = 1'b0;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l176_1) begin
      sram_1_ports_cmd_payload_wen = 16'h0;
    end else begin
      if(when_ICache_l183_1) begin
        sram_1_ports_cmd_payload_wen = 16'h0;
      end else begin
        if(when_ICache_l190_1) begin
          sram_1_ports_cmd_payload_wen = (_zz_sram_1_ports_cmd_payload_wen <<< _zz_sram_1_ports_cmd_payload_wen_1);
        end else begin
          sram_1_ports_cmd_payload_wen = 16'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l176_1) begin
      sram_1_ports_cmd_payload_wdata = 512'h0;
    end else begin
      if(when_ICache_l183_1) begin
        sram_1_ports_cmd_payload_wdata = 512'h0;
      end else begin
        if(when_ICache_l190_1) begin
          sram_1_ports_cmd_payload_wdata = ({448'h0,next_level_rsp_payload_data} <<< _zz_sram_1_ports_cmd_payload_wdata);
        end else begin
          sram_1_ports_cmd_payload_wdata = 512'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l176_1) begin
      sram_1_ports_cmd_payload_wstrb = 64'h0;
    end else begin
      if(when_ICache_l183_1) begin
        sram_1_ports_cmd_payload_wstrb = 64'h0;
      end else begin
        if(when_ICache_l190_1) begin
          sram_1_ports_cmd_payload_wstrb = ({56'h0,8'hff} <<< _zz_sram_1_ports_cmd_payload_wstrb);
        end else begin
          sram_1_ports_cmd_payload_wstrb = 64'h0;
        end
      end
    end
  end

  assign _zz_206 = zz__zz_sram_1_ports_cmd_payload_wen(1'b0);
  always @(*) _zz_sram_1_ports_cmd_payload_wen = _zz_206;
  assign when_ICache_l183_1 = (next_level_done && (2'b01 == evict_id_miss));
  assign when_ICache_l190_1 = (next_level_rsp_valid && (2'b01 == evict_id_miss));
  assign _zz_86 = ({15'd0,1'b1} <<< flush_cnt_value);
  assign _zz_87 = _zz_86[0];
  assign _zz_88 = _zz_86[1];
  assign _zz_89 = _zz_86[2];
  assign _zz_90 = _zz_86[3];
  assign _zz_91 = _zz_86[4];
  assign _zz_92 = _zz_86[5];
  assign _zz_93 = _zz_86[6];
  assign _zz_94 = _zz_86[7];
  assign _zz_95 = _zz_86[8];
  assign _zz_96 = _zz_86[9];
  assign _zz_97 = _zz_86[10];
  assign _zz_98 = _zz_86[11];
  assign _zz_99 = _zz_86[12];
  assign _zz_100 = _zz_86[13];
  assign _zz_101 = _zz_86[14];
  assign _zz_102 = _zz_86[15];
  assign when_ICache_l212_1 = (is_hit && mru_full);
  assign when_ICache_l219_1 = (is_hit && cache_hit_1);
  assign when_ICache_l222_1 = (next_level_done && (2'b01 == evict_id_miss));
  assign when_ICache_l227_1 = (next_level_done && (2'b01 == evict_id_miss));
  assign when_ICache_l232_1 = (flush || is_miss);
  assign when_ICache_l235_1 = (flush_done || next_level_done);
  assign _zz_103 = ({15'd0,1'b1} <<< cpu_set);
  assign _zz_104 = _zz_103[0];
  assign _zz_105 = _zz_103[1];
  assign _zz_106 = _zz_103[2];
  assign _zz_107 = _zz_103[3];
  assign _zz_108 = _zz_103[4];
  assign _zz_109 = _zz_103[5];
  assign _zz_110 = _zz_103[6];
  assign _zz_111 = _zz_103[7];
  assign _zz_112 = _zz_103[8];
  assign _zz_113 = _zz_103[9];
  assign _zz_114 = _zz_103[10];
  assign _zz_115 = _zz_103[11];
  assign _zz_116 = _zz_103[12];
  assign _zz_117 = _zz_103[13];
  assign _zz_118 = _zz_103[14];
  assign _zz_119 = _zz_103[15];
  assign cache_tag_2 = _zz_cache_tag_2;
  assign cache_hit_2 = ((cache_tag_2 == cpu_tag) && _zz_cache_hit_2);
  assign cache_mru_2 = _zz_cache_mru_2;
  assign _zz_120 = ({15'd0,1'b1} <<< cpu_set_d1);
  assign _zz_121 = _zz_120[0];
  assign _zz_122 = _zz_120[1];
  assign _zz_123 = _zz_120[2];
  assign _zz_124 = _zz_120[3];
  assign _zz_125 = _zz_120[4];
  assign _zz_126 = _zz_120[5];
  assign _zz_127 = _zz_120[6];
  assign _zz_128 = _zz_120[7];
  assign _zz_129 = _zz_120[8];
  assign _zz_130 = _zz_120[9];
  assign _zz_131 = _zz_120[10];
  assign _zz_132 = _zz_120[11];
  assign _zz_133 = _zz_120[12];
  assign _zz_134 = _zz_120[13];
  assign _zz_135 = _zz_120[14];
  assign _zz_136 = _zz_120[15];
  assign cache_invld_d1_2 = (! _zz_cache_invld_d1_2);
  assign cache_lru_d1_2 = (! _zz_cache_lru_d1_2);
  assign cache_victim_2 = (cache_invld_d1_2 && cache_lru_d1_2);
  assign sram_banks_data_2 = sram_2_ports_rsp_payload_data;
  assign sram_banks_valid_2 = sram_2_ports_rsp_valid;
  assign when_ICache_l176_2 = (is_hit && (2'b10 == hit_id));
  always @(*) begin
    if(when_ICache_l176_2) begin
      sram_2_ports_cmd_payload_addr = cpu_bank_addr;
    end else begin
      if(when_ICache_l183_2) begin
        sram_2_ports_cmd_payload_addr = cpu_bank_addr_d1;
      end else begin
        if(when_ICache_l190_2) begin
          sram_2_ports_cmd_payload_addr = next_level_bank_addr;
        end else begin
          sram_2_ports_cmd_payload_addr = 4'b0000;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l176_2) begin
      sram_2_ports_cmd_valid = 1'b1;
    end else begin
      if(when_ICache_l183_2) begin
        sram_2_ports_cmd_valid = 1'b1;
      end else begin
        if(when_ICache_l190_2) begin
          sram_2_ports_cmd_valid = 1'b1;
        end else begin
          sram_2_ports_cmd_valid = 1'b0;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l176_2) begin
      sram_2_ports_cmd_payload_wen = 16'h0;
    end else begin
      if(when_ICache_l183_2) begin
        sram_2_ports_cmd_payload_wen = 16'h0;
      end else begin
        if(when_ICache_l190_2) begin
          sram_2_ports_cmd_payload_wen = (_zz_sram_2_ports_cmd_payload_wen <<< _zz_sram_2_ports_cmd_payload_wen_1);
        end else begin
          sram_2_ports_cmd_payload_wen = 16'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l176_2) begin
      sram_2_ports_cmd_payload_wdata = 512'h0;
    end else begin
      if(when_ICache_l183_2) begin
        sram_2_ports_cmd_payload_wdata = 512'h0;
      end else begin
        if(when_ICache_l190_2) begin
          sram_2_ports_cmd_payload_wdata = ({448'h0,next_level_rsp_payload_data} <<< _zz_sram_2_ports_cmd_payload_wdata);
        end else begin
          sram_2_ports_cmd_payload_wdata = 512'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l176_2) begin
      sram_2_ports_cmd_payload_wstrb = 64'h0;
    end else begin
      if(when_ICache_l183_2) begin
        sram_2_ports_cmd_payload_wstrb = 64'h0;
      end else begin
        if(when_ICache_l190_2) begin
          sram_2_ports_cmd_payload_wstrb = ({56'h0,8'hff} <<< _zz_sram_2_ports_cmd_payload_wstrb);
        end else begin
          sram_2_ports_cmd_payload_wstrb = 64'h0;
        end
      end
    end
  end

  assign _zz_207 = zz__zz_sram_2_ports_cmd_payload_wen(1'b0);
  always @(*) _zz_sram_2_ports_cmd_payload_wen = _zz_207;
  assign when_ICache_l183_2 = (next_level_done && (2'b10 == evict_id_miss));
  assign when_ICache_l190_2 = (next_level_rsp_valid && (2'b10 == evict_id_miss));
  assign _zz_137 = ({15'd0,1'b1} <<< flush_cnt_value);
  assign _zz_138 = _zz_137[0];
  assign _zz_139 = _zz_137[1];
  assign _zz_140 = _zz_137[2];
  assign _zz_141 = _zz_137[3];
  assign _zz_142 = _zz_137[4];
  assign _zz_143 = _zz_137[5];
  assign _zz_144 = _zz_137[6];
  assign _zz_145 = _zz_137[7];
  assign _zz_146 = _zz_137[8];
  assign _zz_147 = _zz_137[9];
  assign _zz_148 = _zz_137[10];
  assign _zz_149 = _zz_137[11];
  assign _zz_150 = _zz_137[12];
  assign _zz_151 = _zz_137[13];
  assign _zz_152 = _zz_137[14];
  assign _zz_153 = _zz_137[15];
  assign when_ICache_l212_2 = (is_hit && mru_full);
  assign when_ICache_l219_2 = (is_hit && cache_hit_2);
  assign when_ICache_l222_2 = (next_level_done && (2'b10 == evict_id_miss));
  assign when_ICache_l227_2 = (next_level_done && (2'b10 == evict_id_miss));
  assign when_ICache_l232_2 = (flush || is_miss);
  assign when_ICache_l235_2 = (flush_done || next_level_done);
  assign _zz_154 = ({15'd0,1'b1} <<< cpu_set);
  assign _zz_155 = _zz_154[0];
  assign _zz_156 = _zz_154[1];
  assign _zz_157 = _zz_154[2];
  assign _zz_158 = _zz_154[3];
  assign _zz_159 = _zz_154[4];
  assign _zz_160 = _zz_154[5];
  assign _zz_161 = _zz_154[6];
  assign _zz_162 = _zz_154[7];
  assign _zz_163 = _zz_154[8];
  assign _zz_164 = _zz_154[9];
  assign _zz_165 = _zz_154[10];
  assign _zz_166 = _zz_154[11];
  assign _zz_167 = _zz_154[12];
  assign _zz_168 = _zz_154[13];
  assign _zz_169 = _zz_154[14];
  assign _zz_170 = _zz_154[15];
  assign cache_tag_3 = _zz_cache_tag_3;
  assign cache_hit_3 = ((cache_tag_3 == cpu_tag) && _zz_cache_hit_3);
  assign cache_mru_3 = _zz_cache_mru_3;
  assign _zz_171 = ({15'd0,1'b1} <<< cpu_set_d1);
  assign _zz_172 = _zz_171[0];
  assign _zz_173 = _zz_171[1];
  assign _zz_174 = _zz_171[2];
  assign _zz_175 = _zz_171[3];
  assign _zz_176 = _zz_171[4];
  assign _zz_177 = _zz_171[5];
  assign _zz_178 = _zz_171[6];
  assign _zz_179 = _zz_171[7];
  assign _zz_180 = _zz_171[8];
  assign _zz_181 = _zz_171[9];
  assign _zz_182 = _zz_171[10];
  assign _zz_183 = _zz_171[11];
  assign _zz_184 = _zz_171[12];
  assign _zz_185 = _zz_171[13];
  assign _zz_186 = _zz_171[14];
  assign _zz_187 = _zz_171[15];
  assign cache_invld_d1_3 = (! _zz_cache_invld_d1_3);
  assign cache_lru_d1_3 = (! _zz_cache_lru_d1_3);
  assign cache_victim_3 = (cache_invld_d1_3 && cache_lru_d1_3);
  assign sram_banks_data_3 = sram_3_ports_rsp_payload_data;
  assign sram_banks_valid_3 = sram_3_ports_rsp_valid;
  assign when_ICache_l176_3 = (is_hit && (2'b11 == hit_id));
  always @(*) begin
    if(when_ICache_l176_3) begin
      sram_3_ports_cmd_payload_addr = cpu_bank_addr;
    end else begin
      if(when_ICache_l183_3) begin
        sram_3_ports_cmd_payload_addr = cpu_bank_addr_d1;
      end else begin
        if(when_ICache_l190_3) begin
          sram_3_ports_cmd_payload_addr = next_level_bank_addr;
        end else begin
          sram_3_ports_cmd_payload_addr = 4'b0000;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l176_3) begin
      sram_3_ports_cmd_valid = 1'b1;
    end else begin
      if(when_ICache_l183_3) begin
        sram_3_ports_cmd_valid = 1'b1;
      end else begin
        if(when_ICache_l190_3) begin
          sram_3_ports_cmd_valid = 1'b1;
        end else begin
          sram_3_ports_cmd_valid = 1'b0;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l176_3) begin
      sram_3_ports_cmd_payload_wen = 16'h0;
    end else begin
      if(when_ICache_l183_3) begin
        sram_3_ports_cmd_payload_wen = 16'h0;
      end else begin
        if(when_ICache_l190_3) begin
          sram_3_ports_cmd_payload_wen = (_zz_sram_3_ports_cmd_payload_wen <<< _zz_sram_3_ports_cmd_payload_wen_1);
        end else begin
          sram_3_ports_cmd_payload_wen = 16'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l176_3) begin
      sram_3_ports_cmd_payload_wdata = 512'h0;
    end else begin
      if(when_ICache_l183_3) begin
        sram_3_ports_cmd_payload_wdata = 512'h0;
      end else begin
        if(when_ICache_l190_3) begin
          sram_3_ports_cmd_payload_wdata = ({448'h0,next_level_rsp_payload_data} <<< _zz_sram_3_ports_cmd_payload_wdata);
        end else begin
          sram_3_ports_cmd_payload_wdata = 512'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l176_3) begin
      sram_3_ports_cmd_payload_wstrb = 64'h0;
    end else begin
      if(when_ICache_l183_3) begin
        sram_3_ports_cmd_payload_wstrb = 64'h0;
      end else begin
        if(when_ICache_l190_3) begin
          sram_3_ports_cmd_payload_wstrb = ({56'h0,8'hff} <<< _zz_sram_3_ports_cmd_payload_wstrb);
        end else begin
          sram_3_ports_cmd_payload_wstrb = 64'h0;
        end
      end
    end
  end

  assign _zz_208 = zz__zz_sram_3_ports_cmd_payload_wen(1'b0);
  always @(*) _zz_sram_3_ports_cmd_payload_wen = _zz_208;
  assign when_ICache_l183_3 = (next_level_done && (2'b11 == evict_id_miss));
  assign when_ICache_l190_3 = (next_level_rsp_valid && (2'b11 == evict_id_miss));
  assign _zz_188 = ({15'd0,1'b1} <<< flush_cnt_value);
  assign _zz_189 = _zz_188[0];
  assign _zz_190 = _zz_188[1];
  assign _zz_191 = _zz_188[2];
  assign _zz_192 = _zz_188[3];
  assign _zz_193 = _zz_188[4];
  assign _zz_194 = _zz_188[5];
  assign _zz_195 = _zz_188[6];
  assign _zz_196 = _zz_188[7];
  assign _zz_197 = _zz_188[8];
  assign _zz_198 = _zz_188[9];
  assign _zz_199 = _zz_188[10];
  assign _zz_200 = _zz_188[11];
  assign _zz_201 = _zz_188[12];
  assign _zz_202 = _zz_188[13];
  assign _zz_203 = _zz_188[14];
  assign _zz_204 = _zz_188[15];
  assign when_ICache_l212_3 = (is_hit && mru_full);
  assign when_ICache_l219_3 = (is_hit && cache_hit_3);
  assign when_ICache_l222_3 = (next_level_done && (2'b11 == evict_id_miss));
  assign when_ICache_l227_3 = (next_level_done && (2'b11 == evict_id_miss));
  assign when_ICache_l232_3 = (flush || is_miss);
  assign when_ICache_l235_3 = (flush_done || next_level_done);
  assign _zz_hit_data = _zz__zz_hit_data;
  assign hit_data = _zz_hit_data_1;
  assign _zz_miss_data = _zz__zz_miss_data;
  assign miss_data = _zz_miss_data_1;
  assign cpu_rsp_payload_data = (is_hit_d1 ? hit_data : miss_data);
  assign cpu_rsp_valid = (is_hit_d1 ? _zz_cpu_rsp_valid : _zz_cpu_rsp_valid_1);
  assign cpu_cmd_ready = cpu_cmd_ready_1;
  assign next_level_cmd_payload_addr = {cpu_addr_d1[63 : 6],6'h0};
  assign next_level_cmd_payload_len = 4'b0111;
  assign next_level_cmd_payload_size = 3'b011;
  assign next_level_cmd_valid = next_level_cmd_valid_1;
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      ways_0_metas_0_vld <= 1'b0;
      ways_0_metas_0_tag <= 54'h0;
      ways_0_metas_0_mru <= 1'b0;
      ways_0_metas_1_vld <= 1'b0;
      ways_0_metas_1_tag <= 54'h0;
      ways_0_metas_1_mru <= 1'b0;
      ways_0_metas_2_vld <= 1'b0;
      ways_0_metas_2_tag <= 54'h0;
      ways_0_metas_2_mru <= 1'b0;
      ways_0_metas_3_vld <= 1'b0;
      ways_0_metas_3_tag <= 54'h0;
      ways_0_metas_3_mru <= 1'b0;
      ways_0_metas_4_vld <= 1'b0;
      ways_0_metas_4_tag <= 54'h0;
      ways_0_metas_4_mru <= 1'b0;
      ways_0_metas_5_vld <= 1'b0;
      ways_0_metas_5_tag <= 54'h0;
      ways_0_metas_5_mru <= 1'b0;
      ways_0_metas_6_vld <= 1'b0;
      ways_0_metas_6_tag <= 54'h0;
      ways_0_metas_6_mru <= 1'b0;
      ways_0_metas_7_vld <= 1'b0;
      ways_0_metas_7_tag <= 54'h0;
      ways_0_metas_7_mru <= 1'b0;
      ways_0_metas_8_vld <= 1'b0;
      ways_0_metas_8_tag <= 54'h0;
      ways_0_metas_8_mru <= 1'b0;
      ways_0_metas_9_vld <= 1'b0;
      ways_0_metas_9_tag <= 54'h0;
      ways_0_metas_9_mru <= 1'b0;
      ways_0_metas_10_vld <= 1'b0;
      ways_0_metas_10_tag <= 54'h0;
      ways_0_metas_10_mru <= 1'b0;
      ways_0_metas_11_vld <= 1'b0;
      ways_0_metas_11_tag <= 54'h0;
      ways_0_metas_11_mru <= 1'b0;
      ways_0_metas_12_vld <= 1'b0;
      ways_0_metas_12_tag <= 54'h0;
      ways_0_metas_12_mru <= 1'b0;
      ways_0_metas_13_vld <= 1'b0;
      ways_0_metas_13_tag <= 54'h0;
      ways_0_metas_13_mru <= 1'b0;
      ways_0_metas_14_vld <= 1'b0;
      ways_0_metas_14_tag <= 54'h0;
      ways_0_metas_14_mru <= 1'b0;
      ways_0_metas_15_vld <= 1'b0;
      ways_0_metas_15_tag <= 54'h0;
      ways_0_metas_15_mru <= 1'b0;
      ways_1_metas_0_vld <= 1'b0;
      ways_1_metas_0_tag <= 54'h0;
      ways_1_metas_0_mru <= 1'b0;
      ways_1_metas_1_vld <= 1'b0;
      ways_1_metas_1_tag <= 54'h0;
      ways_1_metas_1_mru <= 1'b0;
      ways_1_metas_2_vld <= 1'b0;
      ways_1_metas_2_tag <= 54'h0;
      ways_1_metas_2_mru <= 1'b0;
      ways_1_metas_3_vld <= 1'b0;
      ways_1_metas_3_tag <= 54'h0;
      ways_1_metas_3_mru <= 1'b0;
      ways_1_metas_4_vld <= 1'b0;
      ways_1_metas_4_tag <= 54'h0;
      ways_1_metas_4_mru <= 1'b0;
      ways_1_metas_5_vld <= 1'b0;
      ways_1_metas_5_tag <= 54'h0;
      ways_1_metas_5_mru <= 1'b0;
      ways_1_metas_6_vld <= 1'b0;
      ways_1_metas_6_tag <= 54'h0;
      ways_1_metas_6_mru <= 1'b0;
      ways_1_metas_7_vld <= 1'b0;
      ways_1_metas_7_tag <= 54'h0;
      ways_1_metas_7_mru <= 1'b0;
      ways_1_metas_8_vld <= 1'b0;
      ways_1_metas_8_tag <= 54'h0;
      ways_1_metas_8_mru <= 1'b0;
      ways_1_metas_9_vld <= 1'b0;
      ways_1_metas_9_tag <= 54'h0;
      ways_1_metas_9_mru <= 1'b0;
      ways_1_metas_10_vld <= 1'b0;
      ways_1_metas_10_tag <= 54'h0;
      ways_1_metas_10_mru <= 1'b0;
      ways_1_metas_11_vld <= 1'b0;
      ways_1_metas_11_tag <= 54'h0;
      ways_1_metas_11_mru <= 1'b0;
      ways_1_metas_12_vld <= 1'b0;
      ways_1_metas_12_tag <= 54'h0;
      ways_1_metas_12_mru <= 1'b0;
      ways_1_metas_13_vld <= 1'b0;
      ways_1_metas_13_tag <= 54'h0;
      ways_1_metas_13_mru <= 1'b0;
      ways_1_metas_14_vld <= 1'b0;
      ways_1_metas_14_tag <= 54'h0;
      ways_1_metas_14_mru <= 1'b0;
      ways_1_metas_15_vld <= 1'b0;
      ways_1_metas_15_tag <= 54'h0;
      ways_1_metas_15_mru <= 1'b0;
      ways_2_metas_0_vld <= 1'b0;
      ways_2_metas_0_tag <= 54'h0;
      ways_2_metas_0_mru <= 1'b0;
      ways_2_metas_1_vld <= 1'b0;
      ways_2_metas_1_tag <= 54'h0;
      ways_2_metas_1_mru <= 1'b0;
      ways_2_metas_2_vld <= 1'b0;
      ways_2_metas_2_tag <= 54'h0;
      ways_2_metas_2_mru <= 1'b0;
      ways_2_metas_3_vld <= 1'b0;
      ways_2_metas_3_tag <= 54'h0;
      ways_2_metas_3_mru <= 1'b0;
      ways_2_metas_4_vld <= 1'b0;
      ways_2_metas_4_tag <= 54'h0;
      ways_2_metas_4_mru <= 1'b0;
      ways_2_metas_5_vld <= 1'b0;
      ways_2_metas_5_tag <= 54'h0;
      ways_2_metas_5_mru <= 1'b0;
      ways_2_metas_6_vld <= 1'b0;
      ways_2_metas_6_tag <= 54'h0;
      ways_2_metas_6_mru <= 1'b0;
      ways_2_metas_7_vld <= 1'b0;
      ways_2_metas_7_tag <= 54'h0;
      ways_2_metas_7_mru <= 1'b0;
      ways_2_metas_8_vld <= 1'b0;
      ways_2_metas_8_tag <= 54'h0;
      ways_2_metas_8_mru <= 1'b0;
      ways_2_metas_9_vld <= 1'b0;
      ways_2_metas_9_tag <= 54'h0;
      ways_2_metas_9_mru <= 1'b0;
      ways_2_metas_10_vld <= 1'b0;
      ways_2_metas_10_tag <= 54'h0;
      ways_2_metas_10_mru <= 1'b0;
      ways_2_metas_11_vld <= 1'b0;
      ways_2_metas_11_tag <= 54'h0;
      ways_2_metas_11_mru <= 1'b0;
      ways_2_metas_12_vld <= 1'b0;
      ways_2_metas_12_tag <= 54'h0;
      ways_2_metas_12_mru <= 1'b0;
      ways_2_metas_13_vld <= 1'b0;
      ways_2_metas_13_tag <= 54'h0;
      ways_2_metas_13_mru <= 1'b0;
      ways_2_metas_14_vld <= 1'b0;
      ways_2_metas_14_tag <= 54'h0;
      ways_2_metas_14_mru <= 1'b0;
      ways_2_metas_15_vld <= 1'b0;
      ways_2_metas_15_tag <= 54'h0;
      ways_2_metas_15_mru <= 1'b0;
      ways_3_metas_0_vld <= 1'b0;
      ways_3_metas_0_tag <= 54'h0;
      ways_3_metas_0_mru <= 1'b0;
      ways_3_metas_1_vld <= 1'b0;
      ways_3_metas_1_tag <= 54'h0;
      ways_3_metas_1_mru <= 1'b0;
      ways_3_metas_2_vld <= 1'b0;
      ways_3_metas_2_tag <= 54'h0;
      ways_3_metas_2_mru <= 1'b0;
      ways_3_metas_3_vld <= 1'b0;
      ways_3_metas_3_tag <= 54'h0;
      ways_3_metas_3_mru <= 1'b0;
      ways_3_metas_4_vld <= 1'b0;
      ways_3_metas_4_tag <= 54'h0;
      ways_3_metas_4_mru <= 1'b0;
      ways_3_metas_5_vld <= 1'b0;
      ways_3_metas_5_tag <= 54'h0;
      ways_3_metas_5_mru <= 1'b0;
      ways_3_metas_6_vld <= 1'b0;
      ways_3_metas_6_tag <= 54'h0;
      ways_3_metas_6_mru <= 1'b0;
      ways_3_metas_7_vld <= 1'b0;
      ways_3_metas_7_tag <= 54'h0;
      ways_3_metas_7_mru <= 1'b0;
      ways_3_metas_8_vld <= 1'b0;
      ways_3_metas_8_tag <= 54'h0;
      ways_3_metas_8_mru <= 1'b0;
      ways_3_metas_9_vld <= 1'b0;
      ways_3_metas_9_tag <= 54'h0;
      ways_3_metas_9_mru <= 1'b0;
      ways_3_metas_10_vld <= 1'b0;
      ways_3_metas_10_tag <= 54'h0;
      ways_3_metas_10_mru <= 1'b0;
      ways_3_metas_11_vld <= 1'b0;
      ways_3_metas_11_tag <= 54'h0;
      ways_3_metas_11_mru <= 1'b0;
      ways_3_metas_12_vld <= 1'b0;
      ways_3_metas_12_tag <= 54'h0;
      ways_3_metas_12_mru <= 1'b0;
      ways_3_metas_13_vld <= 1'b0;
      ways_3_metas_13_tag <= 54'h0;
      ways_3_metas_13_mru <= 1'b0;
      ways_3_metas_14_vld <= 1'b0;
      ways_3_metas_14_tag <= 54'h0;
      ways_3_metas_14_mru <= 1'b0;
      ways_3_metas_15_vld <= 1'b0;
      ways_3_metas_15_tag <= 54'h0;
      ways_3_metas_15_mru <= 1'b0;
      flush_busy <= 1'b0;
      flush_cnt_value <= 4'b0000;
      cpu_addr_d1 <= 64'h0;
      cpu_cmd_ready_1 <= 1'b1;
      next_level_cmd_valid_1 <= 1'b0;
      next_level_data_cnt_value <= 3'b000;
    end else begin
      flush_cnt_value <= flush_cnt_valueNext;
      if(cpu_cmd_fire_2) begin
        cpu_addr_d1 <= cpu_cmd_payload_addr;
      end
      next_level_data_cnt_value <= next_level_data_cnt_valueNext;
      if(is_miss) begin
        next_level_cmd_valid_1 <= 1'b1;
      end else begin
        next_level_cmd_valid_1 <= 1'b0;
      end
      if(flush) begin
        flush_busy <= 1'b1;
      end else begin
        if(flush_done) begin
          flush_busy <= 1'b0;
        end
      end
      if(flush_busy) begin
        if(_zz_36) begin
          ways_0_metas_0_mru <= 1'b0;
        end
        if(_zz_37) begin
          ways_0_metas_1_mru <= 1'b0;
        end
        if(_zz_38) begin
          ways_0_metas_2_mru <= 1'b0;
        end
        if(_zz_39) begin
          ways_0_metas_3_mru <= 1'b0;
        end
        if(_zz_40) begin
          ways_0_metas_4_mru <= 1'b0;
        end
        if(_zz_41) begin
          ways_0_metas_5_mru <= 1'b0;
        end
        if(_zz_42) begin
          ways_0_metas_6_mru <= 1'b0;
        end
        if(_zz_43) begin
          ways_0_metas_7_mru <= 1'b0;
        end
        if(_zz_44) begin
          ways_0_metas_8_mru <= 1'b0;
        end
        if(_zz_45) begin
          ways_0_metas_9_mru <= 1'b0;
        end
        if(_zz_46) begin
          ways_0_metas_10_mru <= 1'b0;
        end
        if(_zz_47) begin
          ways_0_metas_11_mru <= 1'b0;
        end
        if(_zz_48) begin
          ways_0_metas_12_mru <= 1'b0;
        end
        if(_zz_49) begin
          ways_0_metas_13_mru <= 1'b0;
        end
        if(_zz_50) begin
          ways_0_metas_14_mru <= 1'b0;
        end
        if(_zz_51) begin
          ways_0_metas_15_mru <= 1'b0;
        end
        if(_zz_36) begin
          ways_0_metas_0_vld <= 1'b0;
        end
        if(_zz_37) begin
          ways_0_metas_1_vld <= 1'b0;
        end
        if(_zz_38) begin
          ways_0_metas_2_vld <= 1'b0;
        end
        if(_zz_39) begin
          ways_0_metas_3_vld <= 1'b0;
        end
        if(_zz_40) begin
          ways_0_metas_4_vld <= 1'b0;
        end
        if(_zz_41) begin
          ways_0_metas_5_vld <= 1'b0;
        end
        if(_zz_42) begin
          ways_0_metas_6_vld <= 1'b0;
        end
        if(_zz_43) begin
          ways_0_metas_7_vld <= 1'b0;
        end
        if(_zz_44) begin
          ways_0_metas_8_vld <= 1'b0;
        end
        if(_zz_45) begin
          ways_0_metas_9_vld <= 1'b0;
        end
        if(_zz_46) begin
          ways_0_metas_10_vld <= 1'b0;
        end
        if(_zz_47) begin
          ways_0_metas_11_vld <= 1'b0;
        end
        if(_zz_48) begin
          ways_0_metas_12_vld <= 1'b0;
        end
        if(_zz_49) begin
          ways_0_metas_13_vld <= 1'b0;
        end
        if(_zz_50) begin
          ways_0_metas_14_vld <= 1'b0;
        end
        if(_zz_51) begin
          ways_0_metas_15_vld <= 1'b0;
        end
      end else begin
        if(when_ICache_l212) begin
          if(cache_hit_0) begin
            if(_zz_2) begin
              ways_0_metas_0_mru <= 1'b1;
            end
            if(_zz_3) begin
              ways_0_metas_1_mru <= 1'b1;
            end
            if(_zz_4) begin
              ways_0_metas_2_mru <= 1'b1;
            end
            if(_zz_5) begin
              ways_0_metas_3_mru <= 1'b1;
            end
            if(_zz_6) begin
              ways_0_metas_4_mru <= 1'b1;
            end
            if(_zz_7) begin
              ways_0_metas_5_mru <= 1'b1;
            end
            if(_zz_8) begin
              ways_0_metas_6_mru <= 1'b1;
            end
            if(_zz_9) begin
              ways_0_metas_7_mru <= 1'b1;
            end
            if(_zz_10) begin
              ways_0_metas_8_mru <= 1'b1;
            end
            if(_zz_11) begin
              ways_0_metas_9_mru <= 1'b1;
            end
            if(_zz_12) begin
              ways_0_metas_10_mru <= 1'b1;
            end
            if(_zz_13) begin
              ways_0_metas_11_mru <= 1'b1;
            end
            if(_zz_14) begin
              ways_0_metas_12_mru <= 1'b1;
            end
            if(_zz_15) begin
              ways_0_metas_13_mru <= 1'b1;
            end
            if(_zz_16) begin
              ways_0_metas_14_mru <= 1'b1;
            end
            if(_zz_17) begin
              ways_0_metas_15_mru <= 1'b1;
            end
          end else begin
            if(_zz_2) begin
              ways_0_metas_0_mru <= 1'b0;
            end
            if(_zz_3) begin
              ways_0_metas_1_mru <= 1'b0;
            end
            if(_zz_4) begin
              ways_0_metas_2_mru <= 1'b0;
            end
            if(_zz_5) begin
              ways_0_metas_3_mru <= 1'b0;
            end
            if(_zz_6) begin
              ways_0_metas_4_mru <= 1'b0;
            end
            if(_zz_7) begin
              ways_0_metas_5_mru <= 1'b0;
            end
            if(_zz_8) begin
              ways_0_metas_6_mru <= 1'b0;
            end
            if(_zz_9) begin
              ways_0_metas_7_mru <= 1'b0;
            end
            if(_zz_10) begin
              ways_0_metas_8_mru <= 1'b0;
            end
            if(_zz_11) begin
              ways_0_metas_9_mru <= 1'b0;
            end
            if(_zz_12) begin
              ways_0_metas_10_mru <= 1'b0;
            end
            if(_zz_13) begin
              ways_0_metas_11_mru <= 1'b0;
            end
            if(_zz_14) begin
              ways_0_metas_12_mru <= 1'b0;
            end
            if(_zz_15) begin
              ways_0_metas_13_mru <= 1'b0;
            end
            if(_zz_16) begin
              ways_0_metas_14_mru <= 1'b0;
            end
            if(_zz_17) begin
              ways_0_metas_15_mru <= 1'b0;
            end
          end
        end else begin
          if(when_ICache_l219) begin
            if(_zz_2) begin
              ways_0_metas_0_mru <= 1'b1;
            end
            if(_zz_3) begin
              ways_0_metas_1_mru <= 1'b1;
            end
            if(_zz_4) begin
              ways_0_metas_2_mru <= 1'b1;
            end
            if(_zz_5) begin
              ways_0_metas_3_mru <= 1'b1;
            end
            if(_zz_6) begin
              ways_0_metas_4_mru <= 1'b1;
            end
            if(_zz_7) begin
              ways_0_metas_5_mru <= 1'b1;
            end
            if(_zz_8) begin
              ways_0_metas_6_mru <= 1'b1;
            end
            if(_zz_9) begin
              ways_0_metas_7_mru <= 1'b1;
            end
            if(_zz_10) begin
              ways_0_metas_8_mru <= 1'b1;
            end
            if(_zz_11) begin
              ways_0_metas_9_mru <= 1'b1;
            end
            if(_zz_12) begin
              ways_0_metas_10_mru <= 1'b1;
            end
            if(_zz_13) begin
              ways_0_metas_11_mru <= 1'b1;
            end
            if(_zz_14) begin
              ways_0_metas_12_mru <= 1'b1;
            end
            if(_zz_15) begin
              ways_0_metas_13_mru <= 1'b1;
            end
            if(_zz_16) begin
              ways_0_metas_14_mru <= 1'b1;
            end
            if(_zz_17) begin
              ways_0_metas_15_mru <= 1'b1;
            end
          end else begin
            if(when_ICache_l222) begin
              if(_zz_19) begin
                ways_0_metas_0_vld <= 1'b1;
              end
              if(_zz_20) begin
                ways_0_metas_1_vld <= 1'b1;
              end
              if(_zz_21) begin
                ways_0_metas_2_vld <= 1'b1;
              end
              if(_zz_22) begin
                ways_0_metas_3_vld <= 1'b1;
              end
              if(_zz_23) begin
                ways_0_metas_4_vld <= 1'b1;
              end
              if(_zz_24) begin
                ways_0_metas_5_vld <= 1'b1;
              end
              if(_zz_25) begin
                ways_0_metas_6_vld <= 1'b1;
              end
              if(_zz_26) begin
                ways_0_metas_7_vld <= 1'b1;
              end
              if(_zz_27) begin
                ways_0_metas_8_vld <= 1'b1;
              end
              if(_zz_28) begin
                ways_0_metas_9_vld <= 1'b1;
              end
              if(_zz_29) begin
                ways_0_metas_10_vld <= 1'b1;
              end
              if(_zz_30) begin
                ways_0_metas_11_vld <= 1'b1;
              end
              if(_zz_31) begin
                ways_0_metas_12_vld <= 1'b1;
              end
              if(_zz_32) begin
                ways_0_metas_13_vld <= 1'b1;
              end
              if(_zz_33) begin
                ways_0_metas_14_vld <= 1'b1;
              end
              if(_zz_34) begin
                ways_0_metas_15_vld <= 1'b1;
              end
            end
          end
        end
      end
      if(when_ICache_l227) begin
        if(_zz_19) begin
          ways_0_metas_0_tag <= cpu_tag_d1;
        end
        if(_zz_20) begin
          ways_0_metas_1_tag <= cpu_tag_d1;
        end
        if(_zz_21) begin
          ways_0_metas_2_tag <= cpu_tag_d1;
        end
        if(_zz_22) begin
          ways_0_metas_3_tag <= cpu_tag_d1;
        end
        if(_zz_23) begin
          ways_0_metas_4_tag <= cpu_tag_d1;
        end
        if(_zz_24) begin
          ways_0_metas_5_tag <= cpu_tag_d1;
        end
        if(_zz_25) begin
          ways_0_metas_6_tag <= cpu_tag_d1;
        end
        if(_zz_26) begin
          ways_0_metas_7_tag <= cpu_tag_d1;
        end
        if(_zz_27) begin
          ways_0_metas_8_tag <= cpu_tag_d1;
        end
        if(_zz_28) begin
          ways_0_metas_9_tag <= cpu_tag_d1;
        end
        if(_zz_29) begin
          ways_0_metas_10_tag <= cpu_tag_d1;
        end
        if(_zz_30) begin
          ways_0_metas_11_tag <= cpu_tag_d1;
        end
        if(_zz_31) begin
          ways_0_metas_12_tag <= cpu_tag_d1;
        end
        if(_zz_32) begin
          ways_0_metas_13_tag <= cpu_tag_d1;
        end
        if(_zz_33) begin
          ways_0_metas_14_tag <= cpu_tag_d1;
        end
        if(_zz_34) begin
          ways_0_metas_15_tag <= cpu_tag_d1;
        end
      end
      if(when_ICache_l232) begin
        cpu_cmd_ready_1 <= 1'b0;
      end else begin
        if(when_ICache_l235) begin
          cpu_cmd_ready_1 <= 1'b1;
        end
      end
      if(flush_busy) begin
        if(_zz_87) begin
          ways_1_metas_0_mru <= 1'b0;
        end
        if(_zz_88) begin
          ways_1_metas_1_mru <= 1'b0;
        end
        if(_zz_89) begin
          ways_1_metas_2_mru <= 1'b0;
        end
        if(_zz_90) begin
          ways_1_metas_3_mru <= 1'b0;
        end
        if(_zz_91) begin
          ways_1_metas_4_mru <= 1'b0;
        end
        if(_zz_92) begin
          ways_1_metas_5_mru <= 1'b0;
        end
        if(_zz_93) begin
          ways_1_metas_6_mru <= 1'b0;
        end
        if(_zz_94) begin
          ways_1_metas_7_mru <= 1'b0;
        end
        if(_zz_95) begin
          ways_1_metas_8_mru <= 1'b0;
        end
        if(_zz_96) begin
          ways_1_metas_9_mru <= 1'b0;
        end
        if(_zz_97) begin
          ways_1_metas_10_mru <= 1'b0;
        end
        if(_zz_98) begin
          ways_1_metas_11_mru <= 1'b0;
        end
        if(_zz_99) begin
          ways_1_metas_12_mru <= 1'b0;
        end
        if(_zz_100) begin
          ways_1_metas_13_mru <= 1'b0;
        end
        if(_zz_101) begin
          ways_1_metas_14_mru <= 1'b0;
        end
        if(_zz_102) begin
          ways_1_metas_15_mru <= 1'b0;
        end
        if(_zz_87) begin
          ways_1_metas_0_vld <= 1'b0;
        end
        if(_zz_88) begin
          ways_1_metas_1_vld <= 1'b0;
        end
        if(_zz_89) begin
          ways_1_metas_2_vld <= 1'b0;
        end
        if(_zz_90) begin
          ways_1_metas_3_vld <= 1'b0;
        end
        if(_zz_91) begin
          ways_1_metas_4_vld <= 1'b0;
        end
        if(_zz_92) begin
          ways_1_metas_5_vld <= 1'b0;
        end
        if(_zz_93) begin
          ways_1_metas_6_vld <= 1'b0;
        end
        if(_zz_94) begin
          ways_1_metas_7_vld <= 1'b0;
        end
        if(_zz_95) begin
          ways_1_metas_8_vld <= 1'b0;
        end
        if(_zz_96) begin
          ways_1_metas_9_vld <= 1'b0;
        end
        if(_zz_97) begin
          ways_1_metas_10_vld <= 1'b0;
        end
        if(_zz_98) begin
          ways_1_metas_11_vld <= 1'b0;
        end
        if(_zz_99) begin
          ways_1_metas_12_vld <= 1'b0;
        end
        if(_zz_100) begin
          ways_1_metas_13_vld <= 1'b0;
        end
        if(_zz_101) begin
          ways_1_metas_14_vld <= 1'b0;
        end
        if(_zz_102) begin
          ways_1_metas_15_vld <= 1'b0;
        end
      end else begin
        if(when_ICache_l212_1) begin
          if(cache_hit_1) begin
            if(_zz_53) begin
              ways_1_metas_0_mru <= 1'b1;
            end
            if(_zz_54) begin
              ways_1_metas_1_mru <= 1'b1;
            end
            if(_zz_55) begin
              ways_1_metas_2_mru <= 1'b1;
            end
            if(_zz_56) begin
              ways_1_metas_3_mru <= 1'b1;
            end
            if(_zz_57) begin
              ways_1_metas_4_mru <= 1'b1;
            end
            if(_zz_58) begin
              ways_1_metas_5_mru <= 1'b1;
            end
            if(_zz_59) begin
              ways_1_metas_6_mru <= 1'b1;
            end
            if(_zz_60) begin
              ways_1_metas_7_mru <= 1'b1;
            end
            if(_zz_61) begin
              ways_1_metas_8_mru <= 1'b1;
            end
            if(_zz_62) begin
              ways_1_metas_9_mru <= 1'b1;
            end
            if(_zz_63) begin
              ways_1_metas_10_mru <= 1'b1;
            end
            if(_zz_64) begin
              ways_1_metas_11_mru <= 1'b1;
            end
            if(_zz_65) begin
              ways_1_metas_12_mru <= 1'b1;
            end
            if(_zz_66) begin
              ways_1_metas_13_mru <= 1'b1;
            end
            if(_zz_67) begin
              ways_1_metas_14_mru <= 1'b1;
            end
            if(_zz_68) begin
              ways_1_metas_15_mru <= 1'b1;
            end
          end else begin
            if(_zz_53) begin
              ways_1_metas_0_mru <= 1'b0;
            end
            if(_zz_54) begin
              ways_1_metas_1_mru <= 1'b0;
            end
            if(_zz_55) begin
              ways_1_metas_2_mru <= 1'b0;
            end
            if(_zz_56) begin
              ways_1_metas_3_mru <= 1'b0;
            end
            if(_zz_57) begin
              ways_1_metas_4_mru <= 1'b0;
            end
            if(_zz_58) begin
              ways_1_metas_5_mru <= 1'b0;
            end
            if(_zz_59) begin
              ways_1_metas_6_mru <= 1'b0;
            end
            if(_zz_60) begin
              ways_1_metas_7_mru <= 1'b0;
            end
            if(_zz_61) begin
              ways_1_metas_8_mru <= 1'b0;
            end
            if(_zz_62) begin
              ways_1_metas_9_mru <= 1'b0;
            end
            if(_zz_63) begin
              ways_1_metas_10_mru <= 1'b0;
            end
            if(_zz_64) begin
              ways_1_metas_11_mru <= 1'b0;
            end
            if(_zz_65) begin
              ways_1_metas_12_mru <= 1'b0;
            end
            if(_zz_66) begin
              ways_1_metas_13_mru <= 1'b0;
            end
            if(_zz_67) begin
              ways_1_metas_14_mru <= 1'b0;
            end
            if(_zz_68) begin
              ways_1_metas_15_mru <= 1'b0;
            end
          end
        end else begin
          if(when_ICache_l219_1) begin
            if(_zz_53) begin
              ways_1_metas_0_mru <= 1'b1;
            end
            if(_zz_54) begin
              ways_1_metas_1_mru <= 1'b1;
            end
            if(_zz_55) begin
              ways_1_metas_2_mru <= 1'b1;
            end
            if(_zz_56) begin
              ways_1_metas_3_mru <= 1'b1;
            end
            if(_zz_57) begin
              ways_1_metas_4_mru <= 1'b1;
            end
            if(_zz_58) begin
              ways_1_metas_5_mru <= 1'b1;
            end
            if(_zz_59) begin
              ways_1_metas_6_mru <= 1'b1;
            end
            if(_zz_60) begin
              ways_1_metas_7_mru <= 1'b1;
            end
            if(_zz_61) begin
              ways_1_metas_8_mru <= 1'b1;
            end
            if(_zz_62) begin
              ways_1_metas_9_mru <= 1'b1;
            end
            if(_zz_63) begin
              ways_1_metas_10_mru <= 1'b1;
            end
            if(_zz_64) begin
              ways_1_metas_11_mru <= 1'b1;
            end
            if(_zz_65) begin
              ways_1_metas_12_mru <= 1'b1;
            end
            if(_zz_66) begin
              ways_1_metas_13_mru <= 1'b1;
            end
            if(_zz_67) begin
              ways_1_metas_14_mru <= 1'b1;
            end
            if(_zz_68) begin
              ways_1_metas_15_mru <= 1'b1;
            end
          end else begin
            if(when_ICache_l222_1) begin
              if(_zz_70) begin
                ways_1_metas_0_vld <= 1'b1;
              end
              if(_zz_71) begin
                ways_1_metas_1_vld <= 1'b1;
              end
              if(_zz_72) begin
                ways_1_metas_2_vld <= 1'b1;
              end
              if(_zz_73) begin
                ways_1_metas_3_vld <= 1'b1;
              end
              if(_zz_74) begin
                ways_1_metas_4_vld <= 1'b1;
              end
              if(_zz_75) begin
                ways_1_metas_5_vld <= 1'b1;
              end
              if(_zz_76) begin
                ways_1_metas_6_vld <= 1'b1;
              end
              if(_zz_77) begin
                ways_1_metas_7_vld <= 1'b1;
              end
              if(_zz_78) begin
                ways_1_metas_8_vld <= 1'b1;
              end
              if(_zz_79) begin
                ways_1_metas_9_vld <= 1'b1;
              end
              if(_zz_80) begin
                ways_1_metas_10_vld <= 1'b1;
              end
              if(_zz_81) begin
                ways_1_metas_11_vld <= 1'b1;
              end
              if(_zz_82) begin
                ways_1_metas_12_vld <= 1'b1;
              end
              if(_zz_83) begin
                ways_1_metas_13_vld <= 1'b1;
              end
              if(_zz_84) begin
                ways_1_metas_14_vld <= 1'b1;
              end
              if(_zz_85) begin
                ways_1_metas_15_vld <= 1'b1;
              end
            end
          end
        end
      end
      if(when_ICache_l227_1) begin
        if(_zz_70) begin
          ways_1_metas_0_tag <= cpu_tag_d1;
        end
        if(_zz_71) begin
          ways_1_metas_1_tag <= cpu_tag_d1;
        end
        if(_zz_72) begin
          ways_1_metas_2_tag <= cpu_tag_d1;
        end
        if(_zz_73) begin
          ways_1_metas_3_tag <= cpu_tag_d1;
        end
        if(_zz_74) begin
          ways_1_metas_4_tag <= cpu_tag_d1;
        end
        if(_zz_75) begin
          ways_1_metas_5_tag <= cpu_tag_d1;
        end
        if(_zz_76) begin
          ways_1_metas_6_tag <= cpu_tag_d1;
        end
        if(_zz_77) begin
          ways_1_metas_7_tag <= cpu_tag_d1;
        end
        if(_zz_78) begin
          ways_1_metas_8_tag <= cpu_tag_d1;
        end
        if(_zz_79) begin
          ways_1_metas_9_tag <= cpu_tag_d1;
        end
        if(_zz_80) begin
          ways_1_metas_10_tag <= cpu_tag_d1;
        end
        if(_zz_81) begin
          ways_1_metas_11_tag <= cpu_tag_d1;
        end
        if(_zz_82) begin
          ways_1_metas_12_tag <= cpu_tag_d1;
        end
        if(_zz_83) begin
          ways_1_metas_13_tag <= cpu_tag_d1;
        end
        if(_zz_84) begin
          ways_1_metas_14_tag <= cpu_tag_d1;
        end
        if(_zz_85) begin
          ways_1_metas_15_tag <= cpu_tag_d1;
        end
      end
      if(when_ICache_l232_1) begin
        cpu_cmd_ready_1 <= 1'b0;
      end else begin
        if(when_ICache_l235_1) begin
          cpu_cmd_ready_1 <= 1'b1;
        end
      end
      if(flush_busy) begin
        if(_zz_138) begin
          ways_2_metas_0_mru <= 1'b0;
        end
        if(_zz_139) begin
          ways_2_metas_1_mru <= 1'b0;
        end
        if(_zz_140) begin
          ways_2_metas_2_mru <= 1'b0;
        end
        if(_zz_141) begin
          ways_2_metas_3_mru <= 1'b0;
        end
        if(_zz_142) begin
          ways_2_metas_4_mru <= 1'b0;
        end
        if(_zz_143) begin
          ways_2_metas_5_mru <= 1'b0;
        end
        if(_zz_144) begin
          ways_2_metas_6_mru <= 1'b0;
        end
        if(_zz_145) begin
          ways_2_metas_7_mru <= 1'b0;
        end
        if(_zz_146) begin
          ways_2_metas_8_mru <= 1'b0;
        end
        if(_zz_147) begin
          ways_2_metas_9_mru <= 1'b0;
        end
        if(_zz_148) begin
          ways_2_metas_10_mru <= 1'b0;
        end
        if(_zz_149) begin
          ways_2_metas_11_mru <= 1'b0;
        end
        if(_zz_150) begin
          ways_2_metas_12_mru <= 1'b0;
        end
        if(_zz_151) begin
          ways_2_metas_13_mru <= 1'b0;
        end
        if(_zz_152) begin
          ways_2_metas_14_mru <= 1'b0;
        end
        if(_zz_153) begin
          ways_2_metas_15_mru <= 1'b0;
        end
        if(_zz_138) begin
          ways_2_metas_0_vld <= 1'b0;
        end
        if(_zz_139) begin
          ways_2_metas_1_vld <= 1'b0;
        end
        if(_zz_140) begin
          ways_2_metas_2_vld <= 1'b0;
        end
        if(_zz_141) begin
          ways_2_metas_3_vld <= 1'b0;
        end
        if(_zz_142) begin
          ways_2_metas_4_vld <= 1'b0;
        end
        if(_zz_143) begin
          ways_2_metas_5_vld <= 1'b0;
        end
        if(_zz_144) begin
          ways_2_metas_6_vld <= 1'b0;
        end
        if(_zz_145) begin
          ways_2_metas_7_vld <= 1'b0;
        end
        if(_zz_146) begin
          ways_2_metas_8_vld <= 1'b0;
        end
        if(_zz_147) begin
          ways_2_metas_9_vld <= 1'b0;
        end
        if(_zz_148) begin
          ways_2_metas_10_vld <= 1'b0;
        end
        if(_zz_149) begin
          ways_2_metas_11_vld <= 1'b0;
        end
        if(_zz_150) begin
          ways_2_metas_12_vld <= 1'b0;
        end
        if(_zz_151) begin
          ways_2_metas_13_vld <= 1'b0;
        end
        if(_zz_152) begin
          ways_2_metas_14_vld <= 1'b0;
        end
        if(_zz_153) begin
          ways_2_metas_15_vld <= 1'b0;
        end
      end else begin
        if(when_ICache_l212_2) begin
          if(cache_hit_2) begin
            if(_zz_104) begin
              ways_2_metas_0_mru <= 1'b1;
            end
            if(_zz_105) begin
              ways_2_metas_1_mru <= 1'b1;
            end
            if(_zz_106) begin
              ways_2_metas_2_mru <= 1'b1;
            end
            if(_zz_107) begin
              ways_2_metas_3_mru <= 1'b1;
            end
            if(_zz_108) begin
              ways_2_metas_4_mru <= 1'b1;
            end
            if(_zz_109) begin
              ways_2_metas_5_mru <= 1'b1;
            end
            if(_zz_110) begin
              ways_2_metas_6_mru <= 1'b1;
            end
            if(_zz_111) begin
              ways_2_metas_7_mru <= 1'b1;
            end
            if(_zz_112) begin
              ways_2_metas_8_mru <= 1'b1;
            end
            if(_zz_113) begin
              ways_2_metas_9_mru <= 1'b1;
            end
            if(_zz_114) begin
              ways_2_metas_10_mru <= 1'b1;
            end
            if(_zz_115) begin
              ways_2_metas_11_mru <= 1'b1;
            end
            if(_zz_116) begin
              ways_2_metas_12_mru <= 1'b1;
            end
            if(_zz_117) begin
              ways_2_metas_13_mru <= 1'b1;
            end
            if(_zz_118) begin
              ways_2_metas_14_mru <= 1'b1;
            end
            if(_zz_119) begin
              ways_2_metas_15_mru <= 1'b1;
            end
          end else begin
            if(_zz_104) begin
              ways_2_metas_0_mru <= 1'b0;
            end
            if(_zz_105) begin
              ways_2_metas_1_mru <= 1'b0;
            end
            if(_zz_106) begin
              ways_2_metas_2_mru <= 1'b0;
            end
            if(_zz_107) begin
              ways_2_metas_3_mru <= 1'b0;
            end
            if(_zz_108) begin
              ways_2_metas_4_mru <= 1'b0;
            end
            if(_zz_109) begin
              ways_2_metas_5_mru <= 1'b0;
            end
            if(_zz_110) begin
              ways_2_metas_6_mru <= 1'b0;
            end
            if(_zz_111) begin
              ways_2_metas_7_mru <= 1'b0;
            end
            if(_zz_112) begin
              ways_2_metas_8_mru <= 1'b0;
            end
            if(_zz_113) begin
              ways_2_metas_9_mru <= 1'b0;
            end
            if(_zz_114) begin
              ways_2_metas_10_mru <= 1'b0;
            end
            if(_zz_115) begin
              ways_2_metas_11_mru <= 1'b0;
            end
            if(_zz_116) begin
              ways_2_metas_12_mru <= 1'b0;
            end
            if(_zz_117) begin
              ways_2_metas_13_mru <= 1'b0;
            end
            if(_zz_118) begin
              ways_2_metas_14_mru <= 1'b0;
            end
            if(_zz_119) begin
              ways_2_metas_15_mru <= 1'b0;
            end
          end
        end else begin
          if(when_ICache_l219_2) begin
            if(_zz_104) begin
              ways_2_metas_0_mru <= 1'b1;
            end
            if(_zz_105) begin
              ways_2_metas_1_mru <= 1'b1;
            end
            if(_zz_106) begin
              ways_2_metas_2_mru <= 1'b1;
            end
            if(_zz_107) begin
              ways_2_metas_3_mru <= 1'b1;
            end
            if(_zz_108) begin
              ways_2_metas_4_mru <= 1'b1;
            end
            if(_zz_109) begin
              ways_2_metas_5_mru <= 1'b1;
            end
            if(_zz_110) begin
              ways_2_metas_6_mru <= 1'b1;
            end
            if(_zz_111) begin
              ways_2_metas_7_mru <= 1'b1;
            end
            if(_zz_112) begin
              ways_2_metas_8_mru <= 1'b1;
            end
            if(_zz_113) begin
              ways_2_metas_9_mru <= 1'b1;
            end
            if(_zz_114) begin
              ways_2_metas_10_mru <= 1'b1;
            end
            if(_zz_115) begin
              ways_2_metas_11_mru <= 1'b1;
            end
            if(_zz_116) begin
              ways_2_metas_12_mru <= 1'b1;
            end
            if(_zz_117) begin
              ways_2_metas_13_mru <= 1'b1;
            end
            if(_zz_118) begin
              ways_2_metas_14_mru <= 1'b1;
            end
            if(_zz_119) begin
              ways_2_metas_15_mru <= 1'b1;
            end
          end else begin
            if(when_ICache_l222_2) begin
              if(_zz_121) begin
                ways_2_metas_0_vld <= 1'b1;
              end
              if(_zz_122) begin
                ways_2_metas_1_vld <= 1'b1;
              end
              if(_zz_123) begin
                ways_2_metas_2_vld <= 1'b1;
              end
              if(_zz_124) begin
                ways_2_metas_3_vld <= 1'b1;
              end
              if(_zz_125) begin
                ways_2_metas_4_vld <= 1'b1;
              end
              if(_zz_126) begin
                ways_2_metas_5_vld <= 1'b1;
              end
              if(_zz_127) begin
                ways_2_metas_6_vld <= 1'b1;
              end
              if(_zz_128) begin
                ways_2_metas_7_vld <= 1'b1;
              end
              if(_zz_129) begin
                ways_2_metas_8_vld <= 1'b1;
              end
              if(_zz_130) begin
                ways_2_metas_9_vld <= 1'b1;
              end
              if(_zz_131) begin
                ways_2_metas_10_vld <= 1'b1;
              end
              if(_zz_132) begin
                ways_2_metas_11_vld <= 1'b1;
              end
              if(_zz_133) begin
                ways_2_metas_12_vld <= 1'b1;
              end
              if(_zz_134) begin
                ways_2_metas_13_vld <= 1'b1;
              end
              if(_zz_135) begin
                ways_2_metas_14_vld <= 1'b1;
              end
              if(_zz_136) begin
                ways_2_metas_15_vld <= 1'b1;
              end
            end
          end
        end
      end
      if(when_ICache_l227_2) begin
        if(_zz_121) begin
          ways_2_metas_0_tag <= cpu_tag_d1;
        end
        if(_zz_122) begin
          ways_2_metas_1_tag <= cpu_tag_d1;
        end
        if(_zz_123) begin
          ways_2_metas_2_tag <= cpu_tag_d1;
        end
        if(_zz_124) begin
          ways_2_metas_3_tag <= cpu_tag_d1;
        end
        if(_zz_125) begin
          ways_2_metas_4_tag <= cpu_tag_d1;
        end
        if(_zz_126) begin
          ways_2_metas_5_tag <= cpu_tag_d1;
        end
        if(_zz_127) begin
          ways_2_metas_6_tag <= cpu_tag_d1;
        end
        if(_zz_128) begin
          ways_2_metas_7_tag <= cpu_tag_d1;
        end
        if(_zz_129) begin
          ways_2_metas_8_tag <= cpu_tag_d1;
        end
        if(_zz_130) begin
          ways_2_metas_9_tag <= cpu_tag_d1;
        end
        if(_zz_131) begin
          ways_2_metas_10_tag <= cpu_tag_d1;
        end
        if(_zz_132) begin
          ways_2_metas_11_tag <= cpu_tag_d1;
        end
        if(_zz_133) begin
          ways_2_metas_12_tag <= cpu_tag_d1;
        end
        if(_zz_134) begin
          ways_2_metas_13_tag <= cpu_tag_d1;
        end
        if(_zz_135) begin
          ways_2_metas_14_tag <= cpu_tag_d1;
        end
        if(_zz_136) begin
          ways_2_metas_15_tag <= cpu_tag_d1;
        end
      end
      if(when_ICache_l232_2) begin
        cpu_cmd_ready_1 <= 1'b0;
      end else begin
        if(when_ICache_l235_2) begin
          cpu_cmd_ready_1 <= 1'b1;
        end
      end
      if(flush_busy) begin
        if(_zz_189) begin
          ways_3_metas_0_mru <= 1'b0;
        end
        if(_zz_190) begin
          ways_3_metas_1_mru <= 1'b0;
        end
        if(_zz_191) begin
          ways_3_metas_2_mru <= 1'b0;
        end
        if(_zz_192) begin
          ways_3_metas_3_mru <= 1'b0;
        end
        if(_zz_193) begin
          ways_3_metas_4_mru <= 1'b0;
        end
        if(_zz_194) begin
          ways_3_metas_5_mru <= 1'b0;
        end
        if(_zz_195) begin
          ways_3_metas_6_mru <= 1'b0;
        end
        if(_zz_196) begin
          ways_3_metas_7_mru <= 1'b0;
        end
        if(_zz_197) begin
          ways_3_metas_8_mru <= 1'b0;
        end
        if(_zz_198) begin
          ways_3_metas_9_mru <= 1'b0;
        end
        if(_zz_199) begin
          ways_3_metas_10_mru <= 1'b0;
        end
        if(_zz_200) begin
          ways_3_metas_11_mru <= 1'b0;
        end
        if(_zz_201) begin
          ways_3_metas_12_mru <= 1'b0;
        end
        if(_zz_202) begin
          ways_3_metas_13_mru <= 1'b0;
        end
        if(_zz_203) begin
          ways_3_metas_14_mru <= 1'b0;
        end
        if(_zz_204) begin
          ways_3_metas_15_mru <= 1'b0;
        end
        if(_zz_189) begin
          ways_3_metas_0_vld <= 1'b0;
        end
        if(_zz_190) begin
          ways_3_metas_1_vld <= 1'b0;
        end
        if(_zz_191) begin
          ways_3_metas_2_vld <= 1'b0;
        end
        if(_zz_192) begin
          ways_3_metas_3_vld <= 1'b0;
        end
        if(_zz_193) begin
          ways_3_metas_4_vld <= 1'b0;
        end
        if(_zz_194) begin
          ways_3_metas_5_vld <= 1'b0;
        end
        if(_zz_195) begin
          ways_3_metas_6_vld <= 1'b0;
        end
        if(_zz_196) begin
          ways_3_metas_7_vld <= 1'b0;
        end
        if(_zz_197) begin
          ways_3_metas_8_vld <= 1'b0;
        end
        if(_zz_198) begin
          ways_3_metas_9_vld <= 1'b0;
        end
        if(_zz_199) begin
          ways_3_metas_10_vld <= 1'b0;
        end
        if(_zz_200) begin
          ways_3_metas_11_vld <= 1'b0;
        end
        if(_zz_201) begin
          ways_3_metas_12_vld <= 1'b0;
        end
        if(_zz_202) begin
          ways_3_metas_13_vld <= 1'b0;
        end
        if(_zz_203) begin
          ways_3_metas_14_vld <= 1'b0;
        end
        if(_zz_204) begin
          ways_3_metas_15_vld <= 1'b0;
        end
      end else begin
        if(when_ICache_l212_3) begin
          if(cache_hit_3) begin
            if(_zz_155) begin
              ways_3_metas_0_mru <= 1'b1;
            end
            if(_zz_156) begin
              ways_3_metas_1_mru <= 1'b1;
            end
            if(_zz_157) begin
              ways_3_metas_2_mru <= 1'b1;
            end
            if(_zz_158) begin
              ways_3_metas_3_mru <= 1'b1;
            end
            if(_zz_159) begin
              ways_3_metas_4_mru <= 1'b1;
            end
            if(_zz_160) begin
              ways_3_metas_5_mru <= 1'b1;
            end
            if(_zz_161) begin
              ways_3_metas_6_mru <= 1'b1;
            end
            if(_zz_162) begin
              ways_3_metas_7_mru <= 1'b1;
            end
            if(_zz_163) begin
              ways_3_metas_8_mru <= 1'b1;
            end
            if(_zz_164) begin
              ways_3_metas_9_mru <= 1'b1;
            end
            if(_zz_165) begin
              ways_3_metas_10_mru <= 1'b1;
            end
            if(_zz_166) begin
              ways_3_metas_11_mru <= 1'b1;
            end
            if(_zz_167) begin
              ways_3_metas_12_mru <= 1'b1;
            end
            if(_zz_168) begin
              ways_3_metas_13_mru <= 1'b1;
            end
            if(_zz_169) begin
              ways_3_metas_14_mru <= 1'b1;
            end
            if(_zz_170) begin
              ways_3_metas_15_mru <= 1'b1;
            end
          end else begin
            if(_zz_155) begin
              ways_3_metas_0_mru <= 1'b0;
            end
            if(_zz_156) begin
              ways_3_metas_1_mru <= 1'b0;
            end
            if(_zz_157) begin
              ways_3_metas_2_mru <= 1'b0;
            end
            if(_zz_158) begin
              ways_3_metas_3_mru <= 1'b0;
            end
            if(_zz_159) begin
              ways_3_metas_4_mru <= 1'b0;
            end
            if(_zz_160) begin
              ways_3_metas_5_mru <= 1'b0;
            end
            if(_zz_161) begin
              ways_3_metas_6_mru <= 1'b0;
            end
            if(_zz_162) begin
              ways_3_metas_7_mru <= 1'b0;
            end
            if(_zz_163) begin
              ways_3_metas_8_mru <= 1'b0;
            end
            if(_zz_164) begin
              ways_3_metas_9_mru <= 1'b0;
            end
            if(_zz_165) begin
              ways_3_metas_10_mru <= 1'b0;
            end
            if(_zz_166) begin
              ways_3_metas_11_mru <= 1'b0;
            end
            if(_zz_167) begin
              ways_3_metas_12_mru <= 1'b0;
            end
            if(_zz_168) begin
              ways_3_metas_13_mru <= 1'b0;
            end
            if(_zz_169) begin
              ways_3_metas_14_mru <= 1'b0;
            end
            if(_zz_170) begin
              ways_3_metas_15_mru <= 1'b0;
            end
          end
        end else begin
          if(when_ICache_l219_3) begin
            if(_zz_155) begin
              ways_3_metas_0_mru <= 1'b1;
            end
            if(_zz_156) begin
              ways_3_metas_1_mru <= 1'b1;
            end
            if(_zz_157) begin
              ways_3_metas_2_mru <= 1'b1;
            end
            if(_zz_158) begin
              ways_3_metas_3_mru <= 1'b1;
            end
            if(_zz_159) begin
              ways_3_metas_4_mru <= 1'b1;
            end
            if(_zz_160) begin
              ways_3_metas_5_mru <= 1'b1;
            end
            if(_zz_161) begin
              ways_3_metas_6_mru <= 1'b1;
            end
            if(_zz_162) begin
              ways_3_metas_7_mru <= 1'b1;
            end
            if(_zz_163) begin
              ways_3_metas_8_mru <= 1'b1;
            end
            if(_zz_164) begin
              ways_3_metas_9_mru <= 1'b1;
            end
            if(_zz_165) begin
              ways_3_metas_10_mru <= 1'b1;
            end
            if(_zz_166) begin
              ways_3_metas_11_mru <= 1'b1;
            end
            if(_zz_167) begin
              ways_3_metas_12_mru <= 1'b1;
            end
            if(_zz_168) begin
              ways_3_metas_13_mru <= 1'b1;
            end
            if(_zz_169) begin
              ways_3_metas_14_mru <= 1'b1;
            end
            if(_zz_170) begin
              ways_3_metas_15_mru <= 1'b1;
            end
          end else begin
            if(when_ICache_l222_3) begin
              if(_zz_172) begin
                ways_3_metas_0_vld <= 1'b1;
              end
              if(_zz_173) begin
                ways_3_metas_1_vld <= 1'b1;
              end
              if(_zz_174) begin
                ways_3_metas_2_vld <= 1'b1;
              end
              if(_zz_175) begin
                ways_3_metas_3_vld <= 1'b1;
              end
              if(_zz_176) begin
                ways_3_metas_4_vld <= 1'b1;
              end
              if(_zz_177) begin
                ways_3_metas_5_vld <= 1'b1;
              end
              if(_zz_178) begin
                ways_3_metas_6_vld <= 1'b1;
              end
              if(_zz_179) begin
                ways_3_metas_7_vld <= 1'b1;
              end
              if(_zz_180) begin
                ways_3_metas_8_vld <= 1'b1;
              end
              if(_zz_181) begin
                ways_3_metas_9_vld <= 1'b1;
              end
              if(_zz_182) begin
                ways_3_metas_10_vld <= 1'b1;
              end
              if(_zz_183) begin
                ways_3_metas_11_vld <= 1'b1;
              end
              if(_zz_184) begin
                ways_3_metas_12_vld <= 1'b1;
              end
              if(_zz_185) begin
                ways_3_metas_13_vld <= 1'b1;
              end
              if(_zz_186) begin
                ways_3_metas_14_vld <= 1'b1;
              end
              if(_zz_187) begin
                ways_3_metas_15_vld <= 1'b1;
              end
            end
          end
        end
      end
      if(when_ICache_l227_3) begin
        if(_zz_172) begin
          ways_3_metas_0_tag <= cpu_tag_d1;
        end
        if(_zz_173) begin
          ways_3_metas_1_tag <= cpu_tag_d1;
        end
        if(_zz_174) begin
          ways_3_metas_2_tag <= cpu_tag_d1;
        end
        if(_zz_175) begin
          ways_3_metas_3_tag <= cpu_tag_d1;
        end
        if(_zz_176) begin
          ways_3_metas_4_tag <= cpu_tag_d1;
        end
        if(_zz_177) begin
          ways_3_metas_5_tag <= cpu_tag_d1;
        end
        if(_zz_178) begin
          ways_3_metas_6_tag <= cpu_tag_d1;
        end
        if(_zz_179) begin
          ways_3_metas_7_tag <= cpu_tag_d1;
        end
        if(_zz_180) begin
          ways_3_metas_8_tag <= cpu_tag_d1;
        end
        if(_zz_181) begin
          ways_3_metas_9_tag <= cpu_tag_d1;
        end
        if(_zz_182) begin
          ways_3_metas_10_tag <= cpu_tag_d1;
        end
        if(_zz_183) begin
          ways_3_metas_11_tag <= cpu_tag_d1;
        end
        if(_zz_184) begin
          ways_3_metas_12_tag <= cpu_tag_d1;
        end
        if(_zz_185) begin
          ways_3_metas_13_tag <= cpu_tag_d1;
        end
        if(_zz_186) begin
          ways_3_metas_14_tag <= cpu_tag_d1;
        end
        if(_zz_187) begin
          ways_3_metas_15_tag <= cpu_tag_d1;
        end
      end
      if(when_ICache_l232_3) begin
        cpu_cmd_ready_1 <= 1'b0;
      end else begin
        if(when_ICache_l235_3) begin
          cpu_cmd_ready_1 <= 1'b1;
        end
      end
    end
  end

  always @(posedge io_axiClk) begin
    hit_id_d1 <= hit_id;
    is_hit_d1 <= is_hit;
    if(is_miss) begin
      evict_id_miss <= evict_id;
    end
    next_level_done <= (next_level_rsp_valid && (next_level_data_cnt_value == 3'b111));
  end


endmodule

module Timer (
  input               cen,
  input               wen,
  input      [63:0]   addr,
  input      [63:0]   wdata,
  output reg [63:0]   rdata,
  output              timer_int,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  wire       [63:0]   _zz_mtime;
  reg        [63:0]   mtime;
  reg        [63:0]   mtimecmp;
  wire                when_ExcepPlugin_l277;
  wire                when_ExcepPlugin_l290;
  wire                when_ExcepPlugin_l292;

  assign _zz_mtime = (mtime + 64'h0000000000000001);
  assign when_ExcepPlugin_l277 = (wen && cen);
  assign when_ExcepPlugin_l290 = (addr == 64'h000000000200bff8);
  always @(*) begin
    if(when_ExcepPlugin_l290) begin
      rdata = mtime;
    end else begin
      if(when_ExcepPlugin_l292) begin
        rdata = mtimecmp;
      end else begin
        rdata = 64'h0;
      end
    end
  end

  assign when_ExcepPlugin_l292 = (addr == 64'h0000000002004000);
  assign timer_int = (mtimecmp <= mtime);
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      mtime <= 64'h0;
      mtimecmp <= 64'hffffffffffffffff;
    end else begin
      if(when_ExcepPlugin_l277) begin
        case(addr)
          64'h000000000200bff8 : begin
            mtime <= wdata;
          end
          64'h0000000002004000 : begin
            mtimecmp <= wdata;
          end
          default : begin
          end
        endcase
      end else begin
        mtime <= _zz_mtime;
      end
    end
  end


endmodule

module Clint (
  input      [63:0]   pc,
  input      [63:0]   pc_next,
  input               pc_next_valid,
  input               instruction_valid,
  output reg          csr_ports_mepc_wen,
  output reg [63:0]   csr_ports_mepc_wdata,
  output reg          csr_ports_mcause_wen,
  output reg [63:0]   csr_ports_mcause_wdata,
  output reg          csr_ports_mstatus_wen,
  output reg [63:0]   csr_ports_mstatus_wdata,
  input      [63:0]   csr_ports_mtvec,
  input      [63:0]   csr_ports_mepc,
  input      [63:0]   csr_ports_mstatus,
  input               csr_ports_global_int_en,
  input               csr_ports_mtime_int_en,
  input               csr_ports_mtime_int_pend,
  input               timer_int,
  output reg          int_en,
  output reg [63:0]   int_pc,
  output              int_hold,
  input               ecall,
  input               ebreak,
  input               mret,
  input               io_axiClk,
  input               resetCtrl_axiReset
);
  localparam IntTypeEnum_IDLE = 2'd0;
  localparam IntTypeEnum_EXPT = 2'd1;
  localparam IntTypeEnum_TIME_1 = 2'd2;
  localparam IntTypeEnum_MRET = 2'd3;

  reg        [1:0]    int_state;
  reg        [63:0]   pc_next_d1;
  reg        [63:0]   mepc_wdata;
  reg        [63:0]   mcause_wdata;
  wire                when_ExcepPlugin_l180;
  wire                when_ExcepPlugin_l182;
  wire                when_ExcepPlugin_l191;
  wire                when_ExcepPlugin_l208;
  wire                when_ExcepPlugin_l216;

  assign when_ExcepPlugin_l180 = (ecall || ebreak);
  always @(*) begin
    if(when_ExcepPlugin_l180) begin
      int_state = IntTypeEnum_EXPT;
    end else begin
      if(when_ExcepPlugin_l182) begin
        int_state = IntTypeEnum_TIME_1;
      end else begin
        if(mret) begin
          int_state = IntTypeEnum_MRET;
        end else begin
          int_state = IntTypeEnum_IDLE;
        end
      end
    end
  end

  assign when_ExcepPlugin_l182 = ((csr_ports_global_int_en && csr_ports_mtime_int_en) && timer_int);
  assign when_ExcepPlugin_l191 = (int_state == IntTypeEnum_TIME_1);
  always @(*) begin
    if(when_ExcepPlugin_l191) begin
      if(instruction_valid) begin
        mepc_wdata = pc_next;
      end else begin
        mepc_wdata = pc_next_d1;
      end
    end else begin
      if(instruction_valid) begin
        mepc_wdata = pc;
      end else begin
        mepc_wdata = pc_next_d1;
      end
    end
  end

  assign when_ExcepPlugin_l208 = (int_state == IntTypeEnum_EXPT);
  always @(*) begin
    if(when_ExcepPlugin_l208) begin
      if(ecall) begin
        mcause_wdata = 64'h000000000000000b;
      end else begin
        if(ebreak) begin
          mcause_wdata = 64'h0000000000000003;
        end else begin
          mcause_wdata = 64'h000000000000000a;
        end
      end
    end else begin
      if(when_ExcepPlugin_l216) begin
        mcause_wdata = 64'h8000000000000007;
      end else begin
        mcause_wdata = 64'h0;
      end
    end
  end

  assign when_ExcepPlugin_l216 = (int_state == IntTypeEnum_TIME_1);
  always @(*) begin
    if((int_state == IntTypeEnum_EXPT) || (int_state == IntTypeEnum_TIME_1)) begin
        int_en = 1'b1;
    end else if((int_state == IntTypeEnum_MRET)) begin
        int_en = 1'b1;
    end else begin
        int_en = 1'b0;
    end
  end

  always @(*) begin
    if((int_state == IntTypeEnum_EXPT) || (int_state == IntTypeEnum_TIME_1)) begin
        int_pc = csr_ports_mtvec;
    end else if((int_state == IntTypeEnum_MRET)) begin
        int_pc = csr_ports_mepc;
    end else begin
        int_pc = 64'h0;
    end
  end

  always @(*) begin
    if((int_state == IntTypeEnum_EXPT) || (int_state == IntTypeEnum_TIME_1)) begin
        csr_ports_mepc_wen = 1'b1;
    end else if((int_state == IntTypeEnum_MRET)) begin
        csr_ports_mepc_wen = 1'b0;
    end else begin
        csr_ports_mepc_wen = 1'b0;
    end
  end

  always @(*) begin
    if((int_state == IntTypeEnum_EXPT) || (int_state == IntTypeEnum_TIME_1)) begin
        csr_ports_mcause_wen = 1'b1;
    end else if((int_state == IntTypeEnum_MRET)) begin
        csr_ports_mcause_wen = 1'b0;
    end else begin
        csr_ports_mcause_wen = 1'b0;
    end
  end

  always @(*) begin
    if((int_state == IntTypeEnum_EXPT) || (int_state == IntTypeEnum_TIME_1)) begin
        csr_ports_mstatus_wen = 1'b1;
    end else if((int_state == IntTypeEnum_MRET)) begin
        csr_ports_mstatus_wen = 1'b1;
    end else begin
        csr_ports_mstatus_wen = 1'b0;
    end
  end

  always @(*) begin
    if((int_state == IntTypeEnum_EXPT) || (int_state == IntTypeEnum_TIME_1)) begin
        csr_ports_mepc_wdata = mepc_wdata;
    end else if((int_state == IntTypeEnum_MRET)) begin
        csr_ports_mepc_wdata = 64'h0;
    end else begin
        csr_ports_mepc_wdata = 64'h0;
    end
  end

  always @(*) begin
    if((int_state == IntTypeEnum_EXPT) || (int_state == IntTypeEnum_TIME_1)) begin
        csr_ports_mcause_wdata = mcause_wdata;
    end else if((int_state == IntTypeEnum_MRET)) begin
        csr_ports_mcause_wdata = 64'h0;
    end else begin
        csr_ports_mcause_wdata = 64'h0;
    end
  end

  always @(*) begin
    if((int_state == IntTypeEnum_EXPT) || (int_state == IntTypeEnum_TIME_1)) begin
        csr_ports_mstatus_wdata = {{{{csr_ports_mstatus[63 : 8],csr_ports_mstatus[3]},csr_ports_mstatus[6 : 4]},1'b0},csr_ports_mstatus[2 : 0]};
    end else if((int_state == IntTypeEnum_MRET)) begin
        csr_ports_mstatus_wdata = {{{{csr_ports_mstatus[63 : 8],1'b1},csr_ports_mstatus[6 : 4]},csr_ports_mstatus[7]},csr_ports_mstatus[2 : 0]};
    end else begin
        csr_ports_mstatus_wdata = 64'h0;
    end
  end

  assign int_hold = 1'b0;
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      pc_next_d1 <= 64'h0;
    end else begin
      if(pc_next_valid) begin
        pc_next_d1 <= pc_next;
      end
    end
  end


endmodule

module CsrRegfile (
  input      [11:0]   cpu_ports_waddr,
  input               cpu_ports_wen,
  input      [63:0]   cpu_ports_wdata,
  input      [11:0]   cpu_ports_raddr,
  output reg [63:0]   cpu_ports_rdata,
  input               clint_ports_mepc_wen,
  input      [63:0]   clint_ports_mepc_wdata,
  input               clint_ports_mcause_wen,
  input      [63:0]   clint_ports_mcause_wdata,
  input               clint_ports_mstatus_wen,
  input      [63:0]   clint_ports_mstatus_wdata,
  output     [63:0]   clint_ports_mtvec,
  output     [63:0]   clint_ports_mepc,
  output     [63:0]   clint_ports_mstatus,
  output              clint_ports_global_int_en,
  output              clint_ports_mtime_int_en,
  output              clint_ports_mtime_int_pend,
  input               timer_int,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  wire       [63:0]   _zz_mcycle;
  reg        [63:0]   mstatus;
  reg        [63:0]   mie;
  reg        [63:0]   mtvec;
  reg        [63:0]   mepc;
  reg        [63:0]   mcause;
  reg        [63:0]   mtval;
  reg        [63:0]   mip;
  reg        [63:0]   mcycle;
  reg        [63:0]   mhartid;
  reg        [63:0]   mscratch;
  wire                when_ExcepPlugin_l106;

  assign _zz_mcycle = (mcycle + 64'h0000000000000001);
  assign when_ExcepPlugin_l106 = (cpu_ports_wen && (cpu_ports_raddr == cpu_ports_waddr));
  always @(*) begin
    if(when_ExcepPlugin_l106) begin
      cpu_ports_rdata = cpu_ports_wdata;
    end else begin
      case(cpu_ports_raddr)
        12'h300 : begin
          cpu_ports_rdata = mstatus;
        end
        12'h304 : begin
          cpu_ports_rdata = mie;
        end
        12'h305 : begin
          cpu_ports_rdata = mtvec;
        end
        12'h341 : begin
          cpu_ports_rdata = mepc;
        end
        12'h342 : begin
          cpu_ports_rdata = mcause;
        end
        12'h343 : begin
          cpu_ports_rdata = mtval;
        end
        12'h344 : begin
          cpu_ports_rdata = mip;
        end
        12'hb00 : begin
          cpu_ports_rdata = mcycle;
        end
        12'hf14 : begin
          cpu_ports_rdata = mhartid;
        end
        default : begin
          cpu_ports_rdata = 64'h0;
        end
      endcase
    end
  end

  assign clint_ports_mtvec = mtvec;
  assign clint_ports_mepc = mepc;
  assign clint_ports_mstatus = mstatus;
  assign clint_ports_global_int_en = mstatus[3];
  assign clint_ports_mtime_int_en = mie[7];
  assign clint_ports_mtime_int_pend = mip[7];
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      mstatus <= {51'h0,13'h1880};
      mie <= 64'h0;
      mtvec <= 64'h0;
      mepc <= 64'h0;
      mcause <= 64'h0;
      mtval <= 64'h0;
      mip <= 64'h0;
      mcycle <= 64'h0;
      mhartid <= 64'h0;
      mscratch <= 64'h0;
    end else begin
      mcycle <= _zz_mcycle;
      mip <= {{{{52'h0,1'b0},3'b000},timer_int},7'h0};
      if(cpu_ports_wen) begin
        case(cpu_ports_waddr)
          12'h300 : begin
            mstatus <= {{{{{{{((cpu_ports_wdata[16 : 15] == 2'b11) || (cpu_ports_wdata[14 : 13] == 2'b11)),50'h0},2'b11},3'b000},cpu_ports_wdata[7]},3'b000},cpu_ports_wdata[3]},3'b000};
          end
          12'h304 : begin
            mie <= {{{{{{52'h0,cpu_ports_wdata[11]},3'b000},cpu_ports_wdata[7]},3'b000},cpu_ports_wdata[3]},3'b000};
          end
          12'h305 : begin
            mtvec <= cpu_ports_wdata;
          end
          12'h341 : begin
            mepc <= cpu_ports_wdata;
          end
          12'h342 : begin
            mcause <= cpu_ports_wdata;
          end
          12'h343 : begin
            mtval <= cpu_ports_wdata;
          end
          12'hf14 : begin
            mhartid <= cpu_ports_wdata;
          end
          12'h340 : begin
            mscratch <= cpu_ports_wdata;
          end
          default : begin
          end
        endcase
      end else begin
        if(clint_ports_mepc_wen) begin
          mepc <= clint_ports_mepc_wdata;
        end
        if(clint_ports_mcause_wen) begin
          mcause <= clint_ports_mcause_wdata;
        end
        if(clint_ports_mstatus_wen) begin
          mstatus <= clint_ports_mstatus_wdata;
        end
        mtvec <= {clint_ports_mtvec[63 : 2],2'b00};
      end
    end
  end


endmodule

module RegFileModule (
  output     [63:0]   read_ports_rs1_value,
  output     [63:0]   read_ports_rs2_value,
  input      [4:0]    read_ports_rs1_addr,
  input      [4:0]    read_ports_rs2_addr,
  input               read_ports_rs1_req,
  input               read_ports_rs2_req,
  input      [63:0]   write_ports_rd_value,
  input      [4:0]    write_ports_rd_addr,
  input               write_ports_rd_wen,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  reg        [63:0]   _zz_read_value_1;
  reg        [63:0]   _zz_read_value_2;
  reg        [63:0]   reg_file_0;
  reg        [63:0]   reg_file_1;
  reg        [63:0]   reg_file_2;
  reg        [63:0]   reg_file_3;
  reg        [63:0]   reg_file_4;
  reg        [63:0]   reg_file_5;
  reg        [63:0]   reg_file_6;
  reg        [63:0]   reg_file_7;
  reg        [63:0]   reg_file_8;
  reg        [63:0]   reg_file_9;
  reg        [63:0]   reg_file_10;
  reg        [63:0]   reg_file_11;
  reg        [63:0]   reg_file_12;
  reg        [63:0]   reg_file_13;
  reg        [63:0]   reg_file_14;
  reg        [63:0]   reg_file_15;
  reg        [63:0]   reg_file_16;
  reg        [63:0]   reg_file_17;
  reg        [63:0]   reg_file_18;
  reg        [63:0]   reg_file_19;
  reg        [63:0]   reg_file_20;
  reg        [63:0]   reg_file_21;
  reg        [63:0]   reg_file_22;
  reg        [63:0]   reg_file_23;
  reg        [63:0]   reg_file_24;
  reg        [63:0]   reg_file_25;
  reg        [63:0]   reg_file_26;
  reg        [63:0]   reg_file_27;
  reg        [63:0]   reg_file_28;
  reg        [63:0]   reg_file_29;
  reg        [63:0]   reg_file_30;
  reg        [63:0]   reg_file_31;
  wire       [63:0]   read_value_1;
  wire       [63:0]   read_value_2;
  wire                when_DecodePlugin_l61;
  wire       [31:0]   _zz_1;

  always @(*) begin
    case(read_ports_rs1_addr)
      5'b00000 : _zz_read_value_1 = reg_file_0;
      5'b00001 : _zz_read_value_1 = reg_file_1;
      5'b00010 : _zz_read_value_1 = reg_file_2;
      5'b00011 : _zz_read_value_1 = reg_file_3;
      5'b00100 : _zz_read_value_1 = reg_file_4;
      5'b00101 : _zz_read_value_1 = reg_file_5;
      5'b00110 : _zz_read_value_1 = reg_file_6;
      5'b00111 : _zz_read_value_1 = reg_file_7;
      5'b01000 : _zz_read_value_1 = reg_file_8;
      5'b01001 : _zz_read_value_1 = reg_file_9;
      5'b01010 : _zz_read_value_1 = reg_file_10;
      5'b01011 : _zz_read_value_1 = reg_file_11;
      5'b01100 : _zz_read_value_1 = reg_file_12;
      5'b01101 : _zz_read_value_1 = reg_file_13;
      5'b01110 : _zz_read_value_1 = reg_file_14;
      5'b01111 : _zz_read_value_1 = reg_file_15;
      5'b10000 : _zz_read_value_1 = reg_file_16;
      5'b10001 : _zz_read_value_1 = reg_file_17;
      5'b10010 : _zz_read_value_1 = reg_file_18;
      5'b10011 : _zz_read_value_1 = reg_file_19;
      5'b10100 : _zz_read_value_1 = reg_file_20;
      5'b10101 : _zz_read_value_1 = reg_file_21;
      5'b10110 : _zz_read_value_1 = reg_file_22;
      5'b10111 : _zz_read_value_1 = reg_file_23;
      5'b11000 : _zz_read_value_1 = reg_file_24;
      5'b11001 : _zz_read_value_1 = reg_file_25;
      5'b11010 : _zz_read_value_1 = reg_file_26;
      5'b11011 : _zz_read_value_1 = reg_file_27;
      5'b11100 : _zz_read_value_1 = reg_file_28;
      5'b11101 : _zz_read_value_1 = reg_file_29;
      5'b11110 : _zz_read_value_1 = reg_file_30;
      default : _zz_read_value_1 = reg_file_31;
    endcase
  end

  always @(*) begin
    case(read_ports_rs2_addr)
      5'b00000 : _zz_read_value_2 = reg_file_0;
      5'b00001 : _zz_read_value_2 = reg_file_1;
      5'b00010 : _zz_read_value_2 = reg_file_2;
      5'b00011 : _zz_read_value_2 = reg_file_3;
      5'b00100 : _zz_read_value_2 = reg_file_4;
      5'b00101 : _zz_read_value_2 = reg_file_5;
      5'b00110 : _zz_read_value_2 = reg_file_6;
      5'b00111 : _zz_read_value_2 = reg_file_7;
      5'b01000 : _zz_read_value_2 = reg_file_8;
      5'b01001 : _zz_read_value_2 = reg_file_9;
      5'b01010 : _zz_read_value_2 = reg_file_10;
      5'b01011 : _zz_read_value_2 = reg_file_11;
      5'b01100 : _zz_read_value_2 = reg_file_12;
      5'b01101 : _zz_read_value_2 = reg_file_13;
      5'b01110 : _zz_read_value_2 = reg_file_14;
      5'b01111 : _zz_read_value_2 = reg_file_15;
      5'b10000 : _zz_read_value_2 = reg_file_16;
      5'b10001 : _zz_read_value_2 = reg_file_17;
      5'b10010 : _zz_read_value_2 = reg_file_18;
      5'b10011 : _zz_read_value_2 = reg_file_19;
      5'b10100 : _zz_read_value_2 = reg_file_20;
      5'b10101 : _zz_read_value_2 = reg_file_21;
      5'b10110 : _zz_read_value_2 = reg_file_22;
      5'b10111 : _zz_read_value_2 = reg_file_23;
      5'b11000 : _zz_read_value_2 = reg_file_24;
      5'b11001 : _zz_read_value_2 = reg_file_25;
      5'b11010 : _zz_read_value_2 = reg_file_26;
      5'b11011 : _zz_read_value_2 = reg_file_27;
      5'b11100 : _zz_read_value_2 = reg_file_28;
      5'b11101 : _zz_read_value_2 = reg_file_29;
      5'b11110 : _zz_read_value_2 = reg_file_30;
      default : _zz_read_value_2 = reg_file_31;
    endcase
  end

  assign read_value_1 = _zz_read_value_1;
  assign read_value_2 = _zz_read_value_2;
  assign when_DecodePlugin_l61 = (write_ports_rd_wen && (write_ports_rd_addr != 5'h0));
  assign _zz_1 = ({31'd0,1'b1} <<< write_ports_rd_addr);
  assign read_ports_rs1_value = (((write_ports_rd_wen && ((write_ports_rd_addr == read_ports_rs1_addr) && (write_ports_rd_addr != 5'h0))) && read_ports_rs1_req) ? write_ports_rd_value : read_value_1);
  assign read_ports_rs2_value = (((write_ports_rd_wen && ((write_ports_rd_addr == read_ports_rs2_addr) && (write_ports_rd_addr != 5'h0))) && read_ports_rs2_req) ? write_ports_rd_value : read_value_2);
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      reg_file_0 <= 64'h0;
      reg_file_1 <= 64'h0;
      reg_file_2 <= 64'h0;
      reg_file_3 <= 64'h0;
      reg_file_4 <= 64'h0;
      reg_file_5 <= 64'h0;
      reg_file_6 <= 64'h0;
      reg_file_7 <= 64'h0;
      reg_file_8 <= 64'h0;
      reg_file_9 <= 64'h0;
      reg_file_10 <= 64'h0;
      reg_file_11 <= 64'h0;
      reg_file_12 <= 64'h0;
      reg_file_13 <= 64'h0;
      reg_file_14 <= 64'h0;
      reg_file_15 <= 64'h0;
      reg_file_16 <= 64'h0;
      reg_file_17 <= 64'h0;
      reg_file_18 <= 64'h0;
      reg_file_19 <= 64'h0;
      reg_file_20 <= 64'h0;
      reg_file_21 <= 64'h0;
      reg_file_22 <= 64'h0;
      reg_file_23 <= 64'h0;
      reg_file_24 <= 64'h0;
      reg_file_25 <= 64'h0;
      reg_file_26 <= 64'h0;
      reg_file_27 <= 64'h0;
      reg_file_28 <= 64'h0;
      reg_file_29 <= 64'h0;
      reg_file_30 <= 64'h0;
      reg_file_31 <= 64'h0;
    end else begin
      if(when_DecodePlugin_l61) begin
        if(_zz_1[0]) begin
          reg_file_0 <= write_ports_rd_value;
        end
        if(_zz_1[1]) begin
          reg_file_1 <= write_ports_rd_value;
        end
        if(_zz_1[2]) begin
          reg_file_2 <= write_ports_rd_value;
        end
        if(_zz_1[3]) begin
          reg_file_3 <= write_ports_rd_value;
        end
        if(_zz_1[4]) begin
          reg_file_4 <= write_ports_rd_value;
        end
        if(_zz_1[5]) begin
          reg_file_5 <= write_ports_rd_value;
        end
        if(_zz_1[6]) begin
          reg_file_6 <= write_ports_rd_value;
        end
        if(_zz_1[7]) begin
          reg_file_7 <= write_ports_rd_value;
        end
        if(_zz_1[8]) begin
          reg_file_8 <= write_ports_rd_value;
        end
        if(_zz_1[9]) begin
          reg_file_9 <= write_ports_rd_value;
        end
        if(_zz_1[10]) begin
          reg_file_10 <= write_ports_rd_value;
        end
        if(_zz_1[11]) begin
          reg_file_11 <= write_ports_rd_value;
        end
        if(_zz_1[12]) begin
          reg_file_12 <= write_ports_rd_value;
        end
        if(_zz_1[13]) begin
          reg_file_13 <= write_ports_rd_value;
        end
        if(_zz_1[14]) begin
          reg_file_14 <= write_ports_rd_value;
        end
        if(_zz_1[15]) begin
          reg_file_15 <= write_ports_rd_value;
        end
        if(_zz_1[16]) begin
          reg_file_16 <= write_ports_rd_value;
        end
        if(_zz_1[17]) begin
          reg_file_17 <= write_ports_rd_value;
        end
        if(_zz_1[18]) begin
          reg_file_18 <= write_ports_rd_value;
        end
        if(_zz_1[19]) begin
          reg_file_19 <= write_ports_rd_value;
        end
        if(_zz_1[20]) begin
          reg_file_20 <= write_ports_rd_value;
        end
        if(_zz_1[21]) begin
          reg_file_21 <= write_ports_rd_value;
        end
        if(_zz_1[22]) begin
          reg_file_22 <= write_ports_rd_value;
        end
        if(_zz_1[23]) begin
          reg_file_23 <= write_ports_rd_value;
        end
        if(_zz_1[24]) begin
          reg_file_24 <= write_ports_rd_value;
        end
        if(_zz_1[25]) begin
          reg_file_25 <= write_ports_rd_value;
        end
        if(_zz_1[26]) begin
          reg_file_26 <= write_ports_rd_value;
        end
        if(_zz_1[27]) begin
          reg_file_27 <= write_ports_rd_value;
        end
        if(_zz_1[28]) begin
          reg_file_28 <= write_ports_rd_value;
        end
        if(_zz_1[29]) begin
          reg_file_29 <= write_ports_rd_value;
        end
        if(_zz_1[30]) begin
          reg_file_30 <= write_ports_rd_value;
        end
        if(_zz_1[31]) begin
          reg_file_31 <= write_ports_rd_value;
        end
      end
    end
  end


endmodule

module gshare_predictor (
  input      [63:0]   predict_pc,
  input               predict_valid,
  output              predict_taken,
  output     [4:0]    predict_history,
  output     [63:0]   predict_pc_next,
  input               train_valid,
  input               train_taken,
  input               train_mispredicted,
  input      [4:0]    train_history,
  input      [63:0]   train_pc,
  input      [63:0]   train_pc_next,
  input               train_is_call,
  input               train_is_ret,
  input               train_is_jmp,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  reg        [1:0]    _zz_GSHARE_pht_predict_taken;
  reg        [1:0]    _zz_switch_Predictor_l38;
  wire       [3:0]    _zz_BTB_btb_alloc_index_valueNext;
  wire       [0:0]    _zz_BTB_btb_alloc_index_valueNext_1;
  wire       [0:0]    _zz_BTB_btb_is_hit;
  wire       [4:0]    _zz_BTB_btb_is_hit_1;
  wire       [0:0]    _zz_BTB_btb_is_miss;
  wire       [4:0]    _zz_BTB_btb_is_miss_1;
  reg        [63:0]   _zz_RAS_ras_predict_pc;
  wire       [63:0]   _zz_predict_pc_next;
  reg        [4:0]    GSHARE_global_branch_history;
  reg        [1:0]    GSHARE_PHT_0;
  reg        [1:0]    GSHARE_PHT_1;
  reg        [1:0]    GSHARE_PHT_2;
  reg        [1:0]    GSHARE_PHT_3;
  reg        [1:0]    GSHARE_PHT_4;
  reg        [1:0]    GSHARE_PHT_5;
  reg        [1:0]    GSHARE_PHT_6;
  reg        [1:0]    GSHARE_PHT_7;
  reg        [1:0]    GSHARE_PHT_8;
  reg        [1:0]    GSHARE_PHT_9;
  reg        [1:0]    GSHARE_PHT_10;
  reg        [1:0]    GSHARE_PHT_11;
  reg        [1:0]    GSHARE_PHT_12;
  reg        [1:0]    GSHARE_PHT_13;
  reg        [1:0]    GSHARE_PHT_14;
  reg        [1:0]    GSHARE_PHT_15;
  reg        [1:0]    GSHARE_PHT_16;
  reg        [1:0]    GSHARE_PHT_17;
  reg        [1:0]    GSHARE_PHT_18;
  reg        [1:0]    GSHARE_PHT_19;
  reg        [1:0]    GSHARE_PHT_20;
  reg        [1:0]    GSHARE_PHT_21;
  reg        [1:0]    GSHARE_PHT_22;
  reg        [1:0]    GSHARE_PHT_23;
  reg        [1:0]    GSHARE_PHT_24;
  reg        [1:0]    GSHARE_PHT_25;
  reg        [1:0]    GSHARE_PHT_26;
  reg        [1:0]    GSHARE_PHT_27;
  reg        [1:0]    GSHARE_PHT_28;
  reg        [1:0]    GSHARE_PHT_29;
  reg        [1:0]    GSHARE_PHT_30;
  reg        [1:0]    GSHARE_PHT_31;
  wire       [4:0]    GSHARE_predict_index;
  wire       [4:0]    GSHARE_train_index;
  wire                GSHARE_pht_predict_taken;
  wire       [1:0]    switch_Predictor_l38;
  wire       [31:0]   _zz_1;
  wire                _zz_2;
  wire                _zz_3;
  wire                _zz_4;
  wire                _zz_5;
  wire                _zz_6;
  wire                _zz_7;
  wire                _zz_8;
  wire                _zz_9;
  wire                _zz_10;
  wire                _zz_11;
  wire                _zz_12;
  wire                _zz_13;
  wire                _zz_14;
  wire                _zz_15;
  wire                _zz_16;
  wire                _zz_17;
  wire                _zz_18;
  wire                _zz_19;
  wire                _zz_20;
  wire                _zz_21;
  wire                _zz_22;
  wire                _zz_23;
  wire                _zz_24;
  wire                _zz_25;
  wire                _zz_26;
  wire                _zz_27;
  wire                _zz_28;
  wire                _zz_29;
  wire                _zz_30;
  wire                _zz_31;
  wire                _zz_32;
  wire                _zz_33;
  wire                when_Predictor_l61;
  wire                when_Predictor_l70;
  reg        [15:0]   BTB_valid;
  reg        [63:0]   BTB_source_pc_0;
  reg        [63:0]   BTB_source_pc_1;
  reg        [63:0]   BTB_source_pc_2;
  reg        [63:0]   BTB_source_pc_3;
  reg        [63:0]   BTB_source_pc_4;
  reg        [63:0]   BTB_source_pc_5;
  reg        [63:0]   BTB_source_pc_6;
  reg        [63:0]   BTB_source_pc_7;
  reg        [63:0]   BTB_source_pc_8;
  reg        [63:0]   BTB_source_pc_9;
  reg        [63:0]   BTB_source_pc_10;
  reg        [63:0]   BTB_source_pc_11;
  reg        [63:0]   BTB_source_pc_12;
  reg        [63:0]   BTB_source_pc_13;
  reg        [63:0]   BTB_source_pc_14;
  reg        [63:0]   BTB_source_pc_15;
  reg        [15:0]   BTB_call;
  reg        [15:0]   BTB_ret;
  reg        [15:0]   BTB_jmp;
  reg        [63:0]   BTB_target_pc_0;
  reg        [63:0]   BTB_target_pc_1;
  reg        [63:0]   BTB_target_pc_2;
  reg        [63:0]   BTB_target_pc_3;
  reg        [63:0]   BTB_target_pc_4;
  reg        [63:0]   BTB_target_pc_5;
  reg        [63:0]   BTB_target_pc_6;
  reg        [63:0]   BTB_target_pc_7;
  reg        [63:0]   BTB_target_pc_8;
  reg        [63:0]   BTB_target_pc_9;
  reg        [63:0]   BTB_target_pc_10;
  reg        [63:0]   BTB_target_pc_11;
  reg        [63:0]   BTB_target_pc_12;
  reg        [63:0]   BTB_target_pc_13;
  reg        [63:0]   BTB_target_pc_14;
  reg        [63:0]   BTB_target_pc_15;
  reg                 BTB_is_matched;
  reg                 BTB_is_call;
  reg                 BTB_is_ret;
  reg                 BTB_is_jmp;
  reg        [63:0]   BTB_target_pc_read;
  wire                when_Predictor_l95;
  wire                when_Predictor_l95_1;
  wire                when_Predictor_l95_2;
  wire                when_Predictor_l95_3;
  wire                when_Predictor_l95_4;
  wire                when_Predictor_l95_5;
  wire                when_Predictor_l95_6;
  wire                when_Predictor_l95_7;
  wire                when_Predictor_l95_8;
  wire                when_Predictor_l95_9;
  wire                when_Predictor_l95_10;
  wire                when_Predictor_l95_11;
  wire                when_Predictor_l95_12;
  wire                when_Predictor_l95_13;
  wire                when_Predictor_l95_14;
  wire                when_Predictor_l95_15;
  wire       [3:0]    BTB_btb_write_index;
  reg                 BTB_btb_alloc_index_willIncrement;
  reg                 BTB_btb_alloc_index_willClear;
  reg        [3:0]    BTB_btb_alloc_index_valueNext;
  reg        [3:0]    BTB_btb_alloc_index_value;
  wire                BTB_btb_alloc_index_willOverflowIfInc;
  wire                BTB_btb_alloc_index_willOverflow;
  reg                 BTB_btb_is_hit_vec_0;
  reg                 BTB_btb_is_hit_vec_1;
  reg                 BTB_btb_is_hit_vec_2;
  reg                 BTB_btb_is_hit_vec_3;
  reg                 BTB_btb_is_hit_vec_4;
  reg                 BTB_btb_is_hit_vec_5;
  reg                 BTB_btb_is_hit_vec_6;
  reg                 BTB_btb_is_hit_vec_7;
  reg                 BTB_btb_is_hit_vec_8;
  reg                 BTB_btb_is_hit_vec_9;
  reg                 BTB_btb_is_hit_vec_10;
  reg                 BTB_btb_is_hit_vec_11;
  reg                 BTB_btb_is_hit_vec_12;
  reg                 BTB_btb_is_hit_vec_13;
  reg                 BTB_btb_is_hit_vec_14;
  reg                 BTB_btb_is_hit_vec_15;
  reg                 BTB_btb_is_miss_vec_0;
  reg                 BTB_btb_is_miss_vec_1;
  reg                 BTB_btb_is_miss_vec_2;
  reg                 BTB_btb_is_miss_vec_3;
  reg                 BTB_btb_is_miss_vec_4;
  reg                 BTB_btb_is_miss_vec_5;
  reg                 BTB_btb_is_miss_vec_6;
  reg                 BTB_btb_is_miss_vec_7;
  reg                 BTB_btb_is_miss_vec_8;
  reg                 BTB_btb_is_miss_vec_9;
  reg                 BTB_btb_is_miss_vec_10;
  reg                 BTB_btb_is_miss_vec_11;
  reg                 BTB_btb_is_miss_vec_12;
  reg                 BTB_btb_is_miss_vec_13;
  reg                 BTB_btb_is_miss_vec_14;
  reg                 BTB_btb_is_miss_vec_15;
  wire                BTB_btb_is_hit;
  wire                BTB_btb_is_miss;
  wire                when_Predictor_l113;
  wire                when_Predictor_l114;
  wire                when_Predictor_l119;
  wire                when_Predictor_l113_1;
  wire                when_Predictor_l114_1;
  wire                when_Predictor_l119_1;
  wire                when_Predictor_l113_2;
  wire                when_Predictor_l114_2;
  wire                when_Predictor_l119_2;
  wire                when_Predictor_l113_3;
  wire                when_Predictor_l114_3;
  wire                when_Predictor_l119_3;
  wire                when_Predictor_l113_4;
  wire                when_Predictor_l114_4;
  wire                when_Predictor_l119_4;
  wire                when_Predictor_l113_5;
  wire                when_Predictor_l114_5;
  wire                when_Predictor_l119_5;
  wire                when_Predictor_l113_6;
  wire                when_Predictor_l114_6;
  wire                when_Predictor_l119_6;
  wire                when_Predictor_l113_7;
  wire                when_Predictor_l114_7;
  wire                when_Predictor_l119_7;
  wire                when_Predictor_l113_8;
  wire                when_Predictor_l114_8;
  wire                when_Predictor_l119_8;
  wire                when_Predictor_l113_9;
  wire                when_Predictor_l114_9;
  wire                when_Predictor_l119_9;
  wire                when_Predictor_l113_10;
  wire                when_Predictor_l114_10;
  wire                when_Predictor_l119_10;
  wire                when_Predictor_l113_11;
  wire                when_Predictor_l114_11;
  wire                when_Predictor_l119_11;
  wire                when_Predictor_l113_12;
  wire                when_Predictor_l114_12;
  wire                when_Predictor_l119_12;
  wire                when_Predictor_l113_13;
  wire                when_Predictor_l114_13;
  wire                when_Predictor_l119_13;
  wire                when_Predictor_l113_14;
  wire                when_Predictor_l114_14;
  wire                when_Predictor_l119_14;
  wire                when_Predictor_l113_15;
  wire                when_Predictor_l114_15;
  wire                when_Predictor_l119_15;
  wire                _zz_BTB_btb_write_index;
  wire                _zz_BTB_btb_write_index_1;
  wire                _zz_BTB_btb_write_index_2;
  wire                _zz_BTB_btb_write_index_3;
  wire       [15:0]   _zz_34;
  wire       [15:0]   _zz_35;
  wire       [15:0]   _zz_36;
  wire       [15:0]   _zz_37;
  reg        [63:0]   RAS_ras_regfile_0;
  reg        [63:0]   RAS_ras_regfile_1;
  reg        [63:0]   RAS_ras_regfile_2;
  reg        [63:0]   RAS_ras_regfile_3;
  reg        [63:0]   RAS_ras_regfile_4;
  reg        [63:0]   RAS_ras_regfile_5;
  reg        [63:0]   RAS_ras_regfile_6;
  reg        [63:0]   RAS_ras_regfile_7;
  reg        [63:0]   RAS_ras_regfile_8;
  reg        [63:0]   RAS_ras_regfile_9;
  reg        [63:0]   RAS_ras_regfile_10;
  reg        [63:0]   RAS_ras_regfile_11;
  reg        [63:0]   RAS_ras_regfile_12;
  reg        [63:0]   RAS_ras_regfile_13;
  reg        [63:0]   RAS_ras_regfile_14;
  reg        [63:0]   RAS_ras_regfile_15;
  reg        [63:0]   RAS_ras_regfile_16;
  reg        [63:0]   RAS_ras_regfile_17;
  reg        [63:0]   RAS_ras_regfile_18;
  reg        [63:0]   RAS_ras_regfile_19;
  reg        [63:0]   RAS_ras_regfile_20;
  reg        [63:0]   RAS_ras_regfile_21;
  reg        [63:0]   RAS_ras_regfile_22;
  reg        [63:0]   RAS_ras_regfile_23;
  reg        [63:0]   RAS_ras_regfile_24;
  reg        [63:0]   RAS_ras_regfile_25;
  reg        [63:0]   RAS_ras_regfile_26;
  reg        [63:0]   RAS_ras_regfile_27;
  reg        [63:0]   RAS_ras_regfile_28;
  reg        [63:0]   RAS_ras_regfile_29;
  reg        [63:0]   RAS_ras_regfile_30;
  reg        [63:0]   RAS_ras_regfile_31;
  reg        [4:0]    RAS_ras_next_index;
  reg        [4:0]    RAS_ras_curr_index;
  reg        [4:0]    RAS_ras_next_index_proven;
  reg        [4:0]    RAS_ras_curr_index_proven;
  wire       [63:0]   RAS_ras_predict_pc;
  wire                RAS_ras_call_matched;
  wire                RAS_ras_ret_matched;
  wire                when_Predictor_l169;
  wire                when_Predictor_l172;
  wire                when_Predictor_l180;
  wire                when_Predictor_l183;
  wire                when_Predictor_l197;
  wire       [31:0]   _zz_38;
  wire                _zz_39;
  wire                _zz_40;
  wire                _zz_41;
  wire                _zz_42;
  wire                _zz_43;
  wire                _zz_44;
  wire                _zz_45;
  wire                _zz_46;
  wire                _zz_47;
  wire                _zz_48;
  wire                _zz_49;
  wire                _zz_50;
  wire                _zz_51;
  wire                _zz_52;
  wire                _zz_53;
  wire                _zz_54;
  wire                _zz_55;
  wire                _zz_56;
  wire                _zz_57;
  wire                _zz_58;
  wire                _zz_59;
  wire                _zz_60;
  wire                _zz_61;
  wire                _zz_62;
  wire                _zz_63;
  wire                _zz_64;
  wire                _zz_65;
  wire                _zz_66;
  wire                _zz_67;
  wire                _zz_68;
  wire                _zz_69;
  wire                _zz_70;
  wire       [63:0]   _zz_RAS_ras_regfile_0;
  wire       [63:0]   _zz_RAS_ras_regfile_0_1;
  wire                when_Predictor_l205;

  assign _zz_BTB_btb_alloc_index_valueNext_1 = BTB_btb_alloc_index_willIncrement;
  assign _zz_BTB_btb_alloc_index_valueNext = {3'd0, _zz_BTB_btb_alloc_index_valueNext_1};
  assign _zz_predict_pc_next = (predict_pc + 64'h0000000000000004);
  assign _zz_BTB_btb_is_hit = BTB_btb_is_hit_vec_5;
  assign _zz_BTB_btb_is_hit_1 = {BTB_btb_is_hit_vec_4,{BTB_btb_is_hit_vec_3,{BTB_btb_is_hit_vec_2,{BTB_btb_is_hit_vec_1,BTB_btb_is_hit_vec_0}}}};
  assign _zz_BTB_btb_is_miss = BTB_btb_is_miss_vec_5;
  assign _zz_BTB_btb_is_miss_1 = {BTB_btb_is_miss_vec_4,{BTB_btb_is_miss_vec_3,{BTB_btb_is_miss_vec_2,{BTB_btb_is_miss_vec_1,BTB_btb_is_miss_vec_0}}}};
  always @(*) begin
    case(GSHARE_predict_index)
      5'b00000 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_0;
      5'b00001 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_1;
      5'b00010 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_2;
      5'b00011 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_3;
      5'b00100 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_4;
      5'b00101 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_5;
      5'b00110 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_6;
      5'b00111 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_7;
      5'b01000 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_8;
      5'b01001 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_9;
      5'b01010 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_10;
      5'b01011 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_11;
      5'b01100 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_12;
      5'b01101 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_13;
      5'b01110 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_14;
      5'b01111 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_15;
      5'b10000 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_16;
      5'b10001 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_17;
      5'b10010 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_18;
      5'b10011 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_19;
      5'b10100 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_20;
      5'b10101 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_21;
      5'b10110 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_22;
      5'b10111 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_23;
      5'b11000 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_24;
      5'b11001 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_25;
      5'b11010 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_26;
      5'b11011 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_27;
      5'b11100 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_28;
      5'b11101 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_29;
      5'b11110 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_30;
      default : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_31;
    endcase
  end

  always @(*) begin
    case(GSHARE_train_index)
      5'b00000 : _zz_switch_Predictor_l38 = GSHARE_PHT_0;
      5'b00001 : _zz_switch_Predictor_l38 = GSHARE_PHT_1;
      5'b00010 : _zz_switch_Predictor_l38 = GSHARE_PHT_2;
      5'b00011 : _zz_switch_Predictor_l38 = GSHARE_PHT_3;
      5'b00100 : _zz_switch_Predictor_l38 = GSHARE_PHT_4;
      5'b00101 : _zz_switch_Predictor_l38 = GSHARE_PHT_5;
      5'b00110 : _zz_switch_Predictor_l38 = GSHARE_PHT_6;
      5'b00111 : _zz_switch_Predictor_l38 = GSHARE_PHT_7;
      5'b01000 : _zz_switch_Predictor_l38 = GSHARE_PHT_8;
      5'b01001 : _zz_switch_Predictor_l38 = GSHARE_PHT_9;
      5'b01010 : _zz_switch_Predictor_l38 = GSHARE_PHT_10;
      5'b01011 : _zz_switch_Predictor_l38 = GSHARE_PHT_11;
      5'b01100 : _zz_switch_Predictor_l38 = GSHARE_PHT_12;
      5'b01101 : _zz_switch_Predictor_l38 = GSHARE_PHT_13;
      5'b01110 : _zz_switch_Predictor_l38 = GSHARE_PHT_14;
      5'b01111 : _zz_switch_Predictor_l38 = GSHARE_PHT_15;
      5'b10000 : _zz_switch_Predictor_l38 = GSHARE_PHT_16;
      5'b10001 : _zz_switch_Predictor_l38 = GSHARE_PHT_17;
      5'b10010 : _zz_switch_Predictor_l38 = GSHARE_PHT_18;
      5'b10011 : _zz_switch_Predictor_l38 = GSHARE_PHT_19;
      5'b10100 : _zz_switch_Predictor_l38 = GSHARE_PHT_20;
      5'b10101 : _zz_switch_Predictor_l38 = GSHARE_PHT_21;
      5'b10110 : _zz_switch_Predictor_l38 = GSHARE_PHT_22;
      5'b10111 : _zz_switch_Predictor_l38 = GSHARE_PHT_23;
      5'b11000 : _zz_switch_Predictor_l38 = GSHARE_PHT_24;
      5'b11001 : _zz_switch_Predictor_l38 = GSHARE_PHT_25;
      5'b11010 : _zz_switch_Predictor_l38 = GSHARE_PHT_26;
      5'b11011 : _zz_switch_Predictor_l38 = GSHARE_PHT_27;
      5'b11100 : _zz_switch_Predictor_l38 = GSHARE_PHT_28;
      5'b11101 : _zz_switch_Predictor_l38 = GSHARE_PHT_29;
      5'b11110 : _zz_switch_Predictor_l38 = GSHARE_PHT_30;
      default : _zz_switch_Predictor_l38 = GSHARE_PHT_31;
    endcase
  end

  always @(*) begin
    case(RAS_ras_curr_index)
      5'b00000 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_0;
      5'b00001 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_1;
      5'b00010 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_2;
      5'b00011 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_3;
      5'b00100 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_4;
      5'b00101 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_5;
      5'b00110 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_6;
      5'b00111 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_7;
      5'b01000 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_8;
      5'b01001 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_9;
      5'b01010 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_10;
      5'b01011 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_11;
      5'b01100 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_12;
      5'b01101 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_13;
      5'b01110 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_14;
      5'b01111 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_15;
      5'b10000 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_16;
      5'b10001 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_17;
      5'b10010 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_18;
      5'b10011 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_19;
      5'b10100 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_20;
      5'b10101 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_21;
      5'b10110 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_22;
      5'b10111 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_23;
      5'b11000 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_24;
      5'b11001 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_25;
      5'b11010 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_26;
      5'b11011 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_27;
      5'b11100 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_28;
      5'b11101 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_29;
      5'b11110 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_30;
      default : _zz_RAS_ras_predict_pc = RAS_ras_regfile_31;
    endcase
  end

  assign GSHARE_predict_index = (predict_pc[6 : 2] ^ GSHARE_global_branch_history);
  assign GSHARE_train_index = (train_pc[6 : 2] ^ train_history);
  assign GSHARE_pht_predict_taken = _zz_GSHARE_pht_predict_taken[1];
  assign switch_Predictor_l38 = _zz_switch_Predictor_l38;
  assign _zz_1 = ({31'd0,1'b1} <<< GSHARE_train_index);
  assign _zz_2 = _zz_1[0];
  assign _zz_3 = _zz_1[1];
  assign _zz_4 = _zz_1[2];
  assign _zz_5 = _zz_1[3];
  assign _zz_6 = _zz_1[4];
  assign _zz_7 = _zz_1[5];
  assign _zz_8 = _zz_1[6];
  assign _zz_9 = _zz_1[7];
  assign _zz_10 = _zz_1[8];
  assign _zz_11 = _zz_1[9];
  assign _zz_12 = _zz_1[10];
  assign _zz_13 = _zz_1[11];
  assign _zz_14 = _zz_1[12];
  assign _zz_15 = _zz_1[13];
  assign _zz_16 = _zz_1[14];
  assign _zz_17 = _zz_1[15];
  assign _zz_18 = _zz_1[16];
  assign _zz_19 = _zz_1[17];
  assign _zz_20 = _zz_1[18];
  assign _zz_21 = _zz_1[19];
  assign _zz_22 = _zz_1[20];
  assign _zz_23 = _zz_1[21];
  assign _zz_24 = _zz_1[22];
  assign _zz_25 = _zz_1[23];
  assign _zz_26 = _zz_1[24];
  assign _zz_27 = _zz_1[25];
  assign _zz_28 = _zz_1[26];
  assign _zz_29 = _zz_1[27];
  assign _zz_30 = _zz_1[28];
  assign _zz_31 = _zz_1[29];
  assign _zz_32 = _zz_1[30];
  assign _zz_33 = _zz_1[31];
  assign when_Predictor_l61 = (! train_taken);
  assign when_Predictor_l70 = (train_valid && train_mispredicted);
  always @(*) begin
    BTB_is_matched = 1'b0;
    if(when_Predictor_l95) begin
      BTB_is_matched = 1'b1;
    end
    if(when_Predictor_l95_1) begin
      BTB_is_matched = 1'b1;
    end
    if(when_Predictor_l95_2) begin
      BTB_is_matched = 1'b1;
    end
    if(when_Predictor_l95_3) begin
      BTB_is_matched = 1'b1;
    end
    if(when_Predictor_l95_4) begin
      BTB_is_matched = 1'b1;
    end
    if(when_Predictor_l95_5) begin
      BTB_is_matched = 1'b1;
    end
    if(when_Predictor_l95_6) begin
      BTB_is_matched = 1'b1;
    end
    if(when_Predictor_l95_7) begin
      BTB_is_matched = 1'b1;
    end
    if(when_Predictor_l95_8) begin
      BTB_is_matched = 1'b1;
    end
    if(when_Predictor_l95_9) begin
      BTB_is_matched = 1'b1;
    end
    if(when_Predictor_l95_10) begin
      BTB_is_matched = 1'b1;
    end
    if(when_Predictor_l95_11) begin
      BTB_is_matched = 1'b1;
    end
    if(when_Predictor_l95_12) begin
      BTB_is_matched = 1'b1;
    end
    if(when_Predictor_l95_13) begin
      BTB_is_matched = 1'b1;
    end
    if(when_Predictor_l95_14) begin
      BTB_is_matched = 1'b1;
    end
    if(when_Predictor_l95_15) begin
      BTB_is_matched = 1'b1;
    end
  end

  always @(*) begin
    BTB_is_call = 1'b0;
    if(when_Predictor_l95) begin
      BTB_is_call = BTB_call[0];
    end
    if(when_Predictor_l95_1) begin
      BTB_is_call = BTB_call[1];
    end
    if(when_Predictor_l95_2) begin
      BTB_is_call = BTB_call[2];
    end
    if(when_Predictor_l95_3) begin
      BTB_is_call = BTB_call[3];
    end
    if(when_Predictor_l95_4) begin
      BTB_is_call = BTB_call[4];
    end
    if(when_Predictor_l95_5) begin
      BTB_is_call = BTB_call[5];
    end
    if(when_Predictor_l95_6) begin
      BTB_is_call = BTB_call[6];
    end
    if(when_Predictor_l95_7) begin
      BTB_is_call = BTB_call[7];
    end
    if(when_Predictor_l95_8) begin
      BTB_is_call = BTB_call[8];
    end
    if(when_Predictor_l95_9) begin
      BTB_is_call = BTB_call[9];
    end
    if(when_Predictor_l95_10) begin
      BTB_is_call = BTB_call[10];
    end
    if(when_Predictor_l95_11) begin
      BTB_is_call = BTB_call[11];
    end
    if(when_Predictor_l95_12) begin
      BTB_is_call = BTB_call[12];
    end
    if(when_Predictor_l95_13) begin
      BTB_is_call = BTB_call[13];
    end
    if(when_Predictor_l95_14) begin
      BTB_is_call = BTB_call[14];
    end
    if(when_Predictor_l95_15) begin
      BTB_is_call = BTB_call[15];
    end
  end

  always @(*) begin
    BTB_is_ret = 1'b0;
    if(when_Predictor_l95) begin
      BTB_is_ret = BTB_ret[0];
    end
    if(when_Predictor_l95_1) begin
      BTB_is_ret = BTB_ret[1];
    end
    if(when_Predictor_l95_2) begin
      BTB_is_ret = BTB_ret[2];
    end
    if(when_Predictor_l95_3) begin
      BTB_is_ret = BTB_ret[3];
    end
    if(when_Predictor_l95_4) begin
      BTB_is_ret = BTB_ret[4];
    end
    if(when_Predictor_l95_5) begin
      BTB_is_ret = BTB_ret[5];
    end
    if(when_Predictor_l95_6) begin
      BTB_is_ret = BTB_ret[6];
    end
    if(when_Predictor_l95_7) begin
      BTB_is_ret = BTB_ret[7];
    end
    if(when_Predictor_l95_8) begin
      BTB_is_ret = BTB_ret[8];
    end
    if(when_Predictor_l95_9) begin
      BTB_is_ret = BTB_ret[9];
    end
    if(when_Predictor_l95_10) begin
      BTB_is_ret = BTB_ret[10];
    end
    if(when_Predictor_l95_11) begin
      BTB_is_ret = BTB_ret[11];
    end
    if(when_Predictor_l95_12) begin
      BTB_is_ret = BTB_ret[12];
    end
    if(when_Predictor_l95_13) begin
      BTB_is_ret = BTB_ret[13];
    end
    if(when_Predictor_l95_14) begin
      BTB_is_ret = BTB_ret[14];
    end
    if(when_Predictor_l95_15) begin
      BTB_is_ret = BTB_ret[15];
    end
  end

  always @(*) begin
    BTB_is_jmp = 1'b0;
    if(when_Predictor_l95) begin
      BTB_is_jmp = BTB_jmp[0];
    end
    if(when_Predictor_l95_1) begin
      BTB_is_jmp = BTB_jmp[1];
    end
    if(when_Predictor_l95_2) begin
      BTB_is_jmp = BTB_jmp[2];
    end
    if(when_Predictor_l95_3) begin
      BTB_is_jmp = BTB_jmp[3];
    end
    if(when_Predictor_l95_4) begin
      BTB_is_jmp = BTB_jmp[4];
    end
    if(when_Predictor_l95_5) begin
      BTB_is_jmp = BTB_jmp[5];
    end
    if(when_Predictor_l95_6) begin
      BTB_is_jmp = BTB_jmp[6];
    end
    if(when_Predictor_l95_7) begin
      BTB_is_jmp = BTB_jmp[7];
    end
    if(when_Predictor_l95_8) begin
      BTB_is_jmp = BTB_jmp[8];
    end
    if(when_Predictor_l95_9) begin
      BTB_is_jmp = BTB_jmp[9];
    end
    if(when_Predictor_l95_10) begin
      BTB_is_jmp = BTB_jmp[10];
    end
    if(when_Predictor_l95_11) begin
      BTB_is_jmp = BTB_jmp[11];
    end
    if(when_Predictor_l95_12) begin
      BTB_is_jmp = BTB_jmp[12];
    end
    if(when_Predictor_l95_13) begin
      BTB_is_jmp = BTB_jmp[13];
    end
    if(when_Predictor_l95_14) begin
      BTB_is_jmp = BTB_jmp[14];
    end
    if(when_Predictor_l95_15) begin
      BTB_is_jmp = BTB_jmp[15];
    end
  end

  always @(*) begin
    BTB_target_pc_read = 64'h0;
    if(when_Predictor_l95) begin
      BTB_target_pc_read = BTB_target_pc_0;
    end
    if(when_Predictor_l95_1) begin
      BTB_target_pc_read = BTB_target_pc_1;
    end
    if(when_Predictor_l95_2) begin
      BTB_target_pc_read = BTB_target_pc_2;
    end
    if(when_Predictor_l95_3) begin
      BTB_target_pc_read = BTB_target_pc_3;
    end
    if(when_Predictor_l95_4) begin
      BTB_target_pc_read = BTB_target_pc_4;
    end
    if(when_Predictor_l95_5) begin
      BTB_target_pc_read = BTB_target_pc_5;
    end
    if(when_Predictor_l95_6) begin
      BTB_target_pc_read = BTB_target_pc_6;
    end
    if(when_Predictor_l95_7) begin
      BTB_target_pc_read = BTB_target_pc_7;
    end
    if(when_Predictor_l95_8) begin
      BTB_target_pc_read = BTB_target_pc_8;
    end
    if(when_Predictor_l95_9) begin
      BTB_target_pc_read = BTB_target_pc_9;
    end
    if(when_Predictor_l95_10) begin
      BTB_target_pc_read = BTB_target_pc_10;
    end
    if(when_Predictor_l95_11) begin
      BTB_target_pc_read = BTB_target_pc_11;
    end
    if(when_Predictor_l95_12) begin
      BTB_target_pc_read = BTB_target_pc_12;
    end
    if(when_Predictor_l95_13) begin
      BTB_target_pc_read = BTB_target_pc_13;
    end
    if(when_Predictor_l95_14) begin
      BTB_target_pc_read = BTB_target_pc_14;
    end
    if(when_Predictor_l95_15) begin
      BTB_target_pc_read = BTB_target_pc_15;
    end
  end

  assign when_Predictor_l95 = ((BTB_source_pc_0 == predict_pc) && BTB_valid[0]);
  assign when_Predictor_l95_1 = ((BTB_source_pc_1 == predict_pc) && BTB_valid[1]);
  assign when_Predictor_l95_2 = ((BTB_source_pc_2 == predict_pc) && BTB_valid[2]);
  assign when_Predictor_l95_3 = ((BTB_source_pc_3 == predict_pc) && BTB_valid[3]);
  assign when_Predictor_l95_4 = ((BTB_source_pc_4 == predict_pc) && BTB_valid[4]);
  assign when_Predictor_l95_5 = ((BTB_source_pc_5 == predict_pc) && BTB_valid[5]);
  assign when_Predictor_l95_6 = ((BTB_source_pc_6 == predict_pc) && BTB_valid[6]);
  assign when_Predictor_l95_7 = ((BTB_source_pc_7 == predict_pc) && BTB_valid[7]);
  assign when_Predictor_l95_8 = ((BTB_source_pc_8 == predict_pc) && BTB_valid[8]);
  assign when_Predictor_l95_9 = ((BTB_source_pc_9 == predict_pc) && BTB_valid[9]);
  assign when_Predictor_l95_10 = ((BTB_source_pc_10 == predict_pc) && BTB_valid[10]);
  assign when_Predictor_l95_11 = ((BTB_source_pc_11 == predict_pc) && BTB_valid[11]);
  assign when_Predictor_l95_12 = ((BTB_source_pc_12 == predict_pc) && BTB_valid[12]);
  assign when_Predictor_l95_13 = ((BTB_source_pc_13 == predict_pc) && BTB_valid[13]);
  assign when_Predictor_l95_14 = ((BTB_source_pc_14 == predict_pc) && BTB_valid[14]);
  assign when_Predictor_l95_15 = ((BTB_source_pc_15 == predict_pc) && BTB_valid[15]);
  always @(*) begin
    BTB_btb_alloc_index_willIncrement = 1'b0;
    if(BTB_btb_is_miss) begin
      if(!BTB_btb_alloc_index_willOverflowIfInc) begin
        BTB_btb_alloc_index_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    BTB_btb_alloc_index_willClear = 1'b0;
    if(BTB_btb_is_miss) begin
      if(BTB_btb_alloc_index_willOverflowIfInc) begin
        BTB_btb_alloc_index_willClear = 1'b1;
      end
    end
  end

  assign BTB_btb_alloc_index_willOverflowIfInc = (BTB_btb_alloc_index_value == 4'b1111);
  assign BTB_btb_alloc_index_willOverflow = (BTB_btb_alloc_index_willOverflowIfInc && BTB_btb_alloc_index_willIncrement);
  always @(*) begin
    BTB_btb_alloc_index_valueNext = (BTB_btb_alloc_index_value + _zz_BTB_btb_alloc_index_valueNext);
    if(BTB_btb_alloc_index_willClear) begin
      BTB_btb_alloc_index_valueNext = 4'b0000;
    end
  end

  assign BTB_btb_is_hit = (|{BTB_btb_is_hit_vec_15,{BTB_btb_is_hit_vec_14,{BTB_btb_is_hit_vec_13,{BTB_btb_is_hit_vec_12,{BTB_btb_is_hit_vec_11,{BTB_btb_is_hit_vec_10,{BTB_btb_is_hit_vec_9,{BTB_btb_is_hit_vec_8,{BTB_btb_is_hit_vec_7,{BTB_btb_is_hit_vec_6,{_zz_BTB_btb_is_hit,_zz_BTB_btb_is_hit_1}}}}}}}}}}});
  assign BTB_btb_is_miss = (|{BTB_btb_is_miss_vec_15,{BTB_btb_is_miss_vec_14,{BTB_btb_is_miss_vec_13,{BTB_btb_is_miss_vec_12,{BTB_btb_is_miss_vec_11,{BTB_btb_is_miss_vec_10,{BTB_btb_is_miss_vec_9,{BTB_btb_is_miss_vec_8,{BTB_btb_is_miss_vec_7,{BTB_btb_is_miss_vec_6,{_zz_BTB_btb_is_miss,_zz_BTB_btb_is_miss_1}}}}}}}}}}});
  assign when_Predictor_l113 = (train_valid && train_taken);
  assign when_Predictor_l114 = ((BTB_source_pc_0 == train_pc) && BTB_valid[0]);
  always @(*) begin
    if(when_Predictor_l113) begin
      if(when_Predictor_l114) begin
        BTB_btb_is_hit_vec_0 = 1'b1;
      end else begin
        BTB_btb_is_hit_vec_0 = 1'b0;
      end
    end else begin
      BTB_btb_is_hit_vec_0 = 1'b0;
    end
  end

  assign when_Predictor_l119 = ((BTB_source_pc_0 != train_pc) || (! BTB_valid[0]));
  always @(*) begin
    if(when_Predictor_l113) begin
      if(when_Predictor_l119) begin
        BTB_btb_is_miss_vec_0 = 1'b1;
      end else begin
        BTB_btb_is_miss_vec_0 = 1'b0;
      end
    end else begin
      BTB_btb_is_miss_vec_0 = 1'b0;
    end
  end

  assign when_Predictor_l113_1 = (train_valid && train_taken);
  assign when_Predictor_l114_1 = ((BTB_source_pc_1 == train_pc) && BTB_valid[1]);
  always @(*) begin
    if(when_Predictor_l113_1) begin
      if(when_Predictor_l114_1) begin
        BTB_btb_is_hit_vec_1 = 1'b1;
      end else begin
        BTB_btb_is_hit_vec_1 = 1'b0;
      end
    end else begin
      BTB_btb_is_hit_vec_1 = 1'b0;
    end
  end

  assign when_Predictor_l119_1 = ((BTB_source_pc_1 != train_pc) || (! BTB_valid[1]));
  always @(*) begin
    if(when_Predictor_l113_1) begin
      if(when_Predictor_l119_1) begin
        BTB_btb_is_miss_vec_1 = 1'b1;
      end else begin
        BTB_btb_is_miss_vec_1 = 1'b0;
      end
    end else begin
      BTB_btb_is_miss_vec_1 = 1'b0;
    end
  end

  assign when_Predictor_l113_2 = (train_valid && train_taken);
  assign when_Predictor_l114_2 = ((BTB_source_pc_2 == train_pc) && BTB_valid[2]);
  always @(*) begin
    if(when_Predictor_l113_2) begin
      if(when_Predictor_l114_2) begin
        BTB_btb_is_hit_vec_2 = 1'b1;
      end else begin
        BTB_btb_is_hit_vec_2 = 1'b0;
      end
    end else begin
      BTB_btb_is_hit_vec_2 = 1'b0;
    end
  end

  assign when_Predictor_l119_2 = ((BTB_source_pc_2 != train_pc) || (! BTB_valid[2]));
  always @(*) begin
    if(when_Predictor_l113_2) begin
      if(when_Predictor_l119_2) begin
        BTB_btb_is_miss_vec_2 = 1'b1;
      end else begin
        BTB_btb_is_miss_vec_2 = 1'b0;
      end
    end else begin
      BTB_btb_is_miss_vec_2 = 1'b0;
    end
  end

  assign when_Predictor_l113_3 = (train_valid && train_taken);
  assign when_Predictor_l114_3 = ((BTB_source_pc_3 == train_pc) && BTB_valid[3]);
  always @(*) begin
    if(when_Predictor_l113_3) begin
      if(when_Predictor_l114_3) begin
        BTB_btb_is_hit_vec_3 = 1'b1;
      end else begin
        BTB_btb_is_hit_vec_3 = 1'b0;
      end
    end else begin
      BTB_btb_is_hit_vec_3 = 1'b0;
    end
  end

  assign when_Predictor_l119_3 = ((BTB_source_pc_3 != train_pc) || (! BTB_valid[3]));
  always @(*) begin
    if(when_Predictor_l113_3) begin
      if(when_Predictor_l119_3) begin
        BTB_btb_is_miss_vec_3 = 1'b1;
      end else begin
        BTB_btb_is_miss_vec_3 = 1'b0;
      end
    end else begin
      BTB_btb_is_miss_vec_3 = 1'b0;
    end
  end

  assign when_Predictor_l113_4 = (train_valid && train_taken);
  assign when_Predictor_l114_4 = ((BTB_source_pc_4 == train_pc) && BTB_valid[4]);
  always @(*) begin
    if(when_Predictor_l113_4) begin
      if(when_Predictor_l114_4) begin
        BTB_btb_is_hit_vec_4 = 1'b1;
      end else begin
        BTB_btb_is_hit_vec_4 = 1'b0;
      end
    end else begin
      BTB_btb_is_hit_vec_4 = 1'b0;
    end
  end

  assign when_Predictor_l119_4 = ((BTB_source_pc_4 != train_pc) || (! BTB_valid[4]));
  always @(*) begin
    if(when_Predictor_l113_4) begin
      if(when_Predictor_l119_4) begin
        BTB_btb_is_miss_vec_4 = 1'b1;
      end else begin
        BTB_btb_is_miss_vec_4 = 1'b0;
      end
    end else begin
      BTB_btb_is_miss_vec_4 = 1'b0;
    end
  end

  assign when_Predictor_l113_5 = (train_valid && train_taken);
  assign when_Predictor_l114_5 = ((BTB_source_pc_5 == train_pc) && BTB_valid[5]);
  always @(*) begin
    if(when_Predictor_l113_5) begin
      if(when_Predictor_l114_5) begin
        BTB_btb_is_hit_vec_5 = 1'b1;
      end else begin
        BTB_btb_is_hit_vec_5 = 1'b0;
      end
    end else begin
      BTB_btb_is_hit_vec_5 = 1'b0;
    end
  end

  assign when_Predictor_l119_5 = ((BTB_source_pc_5 != train_pc) || (! BTB_valid[5]));
  always @(*) begin
    if(when_Predictor_l113_5) begin
      if(when_Predictor_l119_5) begin
        BTB_btb_is_miss_vec_5 = 1'b1;
      end else begin
        BTB_btb_is_miss_vec_5 = 1'b0;
      end
    end else begin
      BTB_btb_is_miss_vec_5 = 1'b0;
    end
  end

  assign when_Predictor_l113_6 = (train_valid && train_taken);
  assign when_Predictor_l114_6 = ((BTB_source_pc_6 == train_pc) && BTB_valid[6]);
  always @(*) begin
    if(when_Predictor_l113_6) begin
      if(when_Predictor_l114_6) begin
        BTB_btb_is_hit_vec_6 = 1'b1;
      end else begin
        BTB_btb_is_hit_vec_6 = 1'b0;
      end
    end else begin
      BTB_btb_is_hit_vec_6 = 1'b0;
    end
  end

  assign when_Predictor_l119_6 = ((BTB_source_pc_6 != train_pc) || (! BTB_valid[6]));
  always @(*) begin
    if(when_Predictor_l113_6) begin
      if(when_Predictor_l119_6) begin
        BTB_btb_is_miss_vec_6 = 1'b1;
      end else begin
        BTB_btb_is_miss_vec_6 = 1'b0;
      end
    end else begin
      BTB_btb_is_miss_vec_6 = 1'b0;
    end
  end

  assign when_Predictor_l113_7 = (train_valid && train_taken);
  assign when_Predictor_l114_7 = ((BTB_source_pc_7 == train_pc) && BTB_valid[7]);
  always @(*) begin
    if(when_Predictor_l113_7) begin
      if(when_Predictor_l114_7) begin
        BTB_btb_is_hit_vec_7 = 1'b1;
      end else begin
        BTB_btb_is_hit_vec_7 = 1'b0;
      end
    end else begin
      BTB_btb_is_hit_vec_7 = 1'b0;
    end
  end

  assign when_Predictor_l119_7 = ((BTB_source_pc_7 != train_pc) || (! BTB_valid[7]));
  always @(*) begin
    if(when_Predictor_l113_7) begin
      if(when_Predictor_l119_7) begin
        BTB_btb_is_miss_vec_7 = 1'b1;
      end else begin
        BTB_btb_is_miss_vec_7 = 1'b0;
      end
    end else begin
      BTB_btb_is_miss_vec_7 = 1'b0;
    end
  end

  assign when_Predictor_l113_8 = (train_valid && train_taken);
  assign when_Predictor_l114_8 = ((BTB_source_pc_8 == train_pc) && BTB_valid[8]);
  always @(*) begin
    if(when_Predictor_l113_8) begin
      if(when_Predictor_l114_8) begin
        BTB_btb_is_hit_vec_8 = 1'b1;
      end else begin
        BTB_btb_is_hit_vec_8 = 1'b0;
      end
    end else begin
      BTB_btb_is_hit_vec_8 = 1'b0;
    end
  end

  assign when_Predictor_l119_8 = ((BTB_source_pc_8 != train_pc) || (! BTB_valid[8]));
  always @(*) begin
    if(when_Predictor_l113_8) begin
      if(when_Predictor_l119_8) begin
        BTB_btb_is_miss_vec_8 = 1'b1;
      end else begin
        BTB_btb_is_miss_vec_8 = 1'b0;
      end
    end else begin
      BTB_btb_is_miss_vec_8 = 1'b0;
    end
  end

  assign when_Predictor_l113_9 = (train_valid && train_taken);
  assign when_Predictor_l114_9 = ((BTB_source_pc_9 == train_pc) && BTB_valid[9]);
  always @(*) begin
    if(when_Predictor_l113_9) begin
      if(when_Predictor_l114_9) begin
        BTB_btb_is_hit_vec_9 = 1'b1;
      end else begin
        BTB_btb_is_hit_vec_9 = 1'b0;
      end
    end else begin
      BTB_btb_is_hit_vec_9 = 1'b0;
    end
  end

  assign when_Predictor_l119_9 = ((BTB_source_pc_9 != train_pc) || (! BTB_valid[9]));
  always @(*) begin
    if(when_Predictor_l113_9) begin
      if(when_Predictor_l119_9) begin
        BTB_btb_is_miss_vec_9 = 1'b1;
      end else begin
        BTB_btb_is_miss_vec_9 = 1'b0;
      end
    end else begin
      BTB_btb_is_miss_vec_9 = 1'b0;
    end
  end

  assign when_Predictor_l113_10 = (train_valid && train_taken);
  assign when_Predictor_l114_10 = ((BTB_source_pc_10 == train_pc) && BTB_valid[10]);
  always @(*) begin
    if(when_Predictor_l113_10) begin
      if(when_Predictor_l114_10) begin
        BTB_btb_is_hit_vec_10 = 1'b1;
      end else begin
        BTB_btb_is_hit_vec_10 = 1'b0;
      end
    end else begin
      BTB_btb_is_hit_vec_10 = 1'b0;
    end
  end

  assign when_Predictor_l119_10 = ((BTB_source_pc_10 != train_pc) || (! BTB_valid[10]));
  always @(*) begin
    if(when_Predictor_l113_10) begin
      if(when_Predictor_l119_10) begin
        BTB_btb_is_miss_vec_10 = 1'b1;
      end else begin
        BTB_btb_is_miss_vec_10 = 1'b0;
      end
    end else begin
      BTB_btb_is_miss_vec_10 = 1'b0;
    end
  end

  assign when_Predictor_l113_11 = (train_valid && train_taken);
  assign when_Predictor_l114_11 = ((BTB_source_pc_11 == train_pc) && BTB_valid[11]);
  always @(*) begin
    if(when_Predictor_l113_11) begin
      if(when_Predictor_l114_11) begin
        BTB_btb_is_hit_vec_11 = 1'b1;
      end else begin
        BTB_btb_is_hit_vec_11 = 1'b0;
      end
    end else begin
      BTB_btb_is_hit_vec_11 = 1'b0;
    end
  end

  assign when_Predictor_l119_11 = ((BTB_source_pc_11 != train_pc) || (! BTB_valid[11]));
  always @(*) begin
    if(when_Predictor_l113_11) begin
      if(when_Predictor_l119_11) begin
        BTB_btb_is_miss_vec_11 = 1'b1;
      end else begin
        BTB_btb_is_miss_vec_11 = 1'b0;
      end
    end else begin
      BTB_btb_is_miss_vec_11 = 1'b0;
    end
  end

  assign when_Predictor_l113_12 = (train_valid && train_taken);
  assign when_Predictor_l114_12 = ((BTB_source_pc_12 == train_pc) && BTB_valid[12]);
  always @(*) begin
    if(when_Predictor_l113_12) begin
      if(when_Predictor_l114_12) begin
        BTB_btb_is_hit_vec_12 = 1'b1;
      end else begin
        BTB_btb_is_hit_vec_12 = 1'b0;
      end
    end else begin
      BTB_btb_is_hit_vec_12 = 1'b0;
    end
  end

  assign when_Predictor_l119_12 = ((BTB_source_pc_12 != train_pc) || (! BTB_valid[12]));
  always @(*) begin
    if(when_Predictor_l113_12) begin
      if(when_Predictor_l119_12) begin
        BTB_btb_is_miss_vec_12 = 1'b1;
      end else begin
        BTB_btb_is_miss_vec_12 = 1'b0;
      end
    end else begin
      BTB_btb_is_miss_vec_12 = 1'b0;
    end
  end

  assign when_Predictor_l113_13 = (train_valid && train_taken);
  assign when_Predictor_l114_13 = ((BTB_source_pc_13 == train_pc) && BTB_valid[13]);
  always @(*) begin
    if(when_Predictor_l113_13) begin
      if(when_Predictor_l114_13) begin
        BTB_btb_is_hit_vec_13 = 1'b1;
      end else begin
        BTB_btb_is_hit_vec_13 = 1'b0;
      end
    end else begin
      BTB_btb_is_hit_vec_13 = 1'b0;
    end
  end

  assign when_Predictor_l119_13 = ((BTB_source_pc_13 != train_pc) || (! BTB_valid[13]));
  always @(*) begin
    if(when_Predictor_l113_13) begin
      if(when_Predictor_l119_13) begin
        BTB_btb_is_miss_vec_13 = 1'b1;
      end else begin
        BTB_btb_is_miss_vec_13 = 1'b0;
      end
    end else begin
      BTB_btb_is_miss_vec_13 = 1'b0;
    end
  end

  assign when_Predictor_l113_14 = (train_valid && train_taken);
  assign when_Predictor_l114_14 = ((BTB_source_pc_14 == train_pc) && BTB_valid[14]);
  always @(*) begin
    if(when_Predictor_l113_14) begin
      if(when_Predictor_l114_14) begin
        BTB_btb_is_hit_vec_14 = 1'b1;
      end else begin
        BTB_btb_is_hit_vec_14 = 1'b0;
      end
    end else begin
      BTB_btb_is_hit_vec_14 = 1'b0;
    end
  end

  assign when_Predictor_l119_14 = ((BTB_source_pc_14 != train_pc) || (! BTB_valid[14]));
  always @(*) begin
    if(when_Predictor_l113_14) begin
      if(when_Predictor_l119_14) begin
        BTB_btb_is_miss_vec_14 = 1'b1;
      end else begin
        BTB_btb_is_miss_vec_14 = 1'b0;
      end
    end else begin
      BTB_btb_is_miss_vec_14 = 1'b0;
    end
  end

  assign when_Predictor_l113_15 = (train_valid && train_taken);
  assign when_Predictor_l114_15 = ((BTB_source_pc_15 == train_pc) && BTB_valid[15]);
  always @(*) begin
    if(when_Predictor_l113_15) begin
      if(when_Predictor_l114_15) begin
        BTB_btb_is_hit_vec_15 = 1'b1;
      end else begin
        BTB_btb_is_hit_vec_15 = 1'b0;
      end
    end else begin
      BTB_btb_is_hit_vec_15 = 1'b0;
    end
  end

  assign when_Predictor_l119_15 = ((BTB_source_pc_15 != train_pc) || (! BTB_valid[15]));
  always @(*) begin
    if(when_Predictor_l113_15) begin
      if(when_Predictor_l119_15) begin
        BTB_btb_is_miss_vec_15 = 1'b1;
      end else begin
        BTB_btb_is_miss_vec_15 = 1'b0;
      end
    end else begin
      BTB_btb_is_miss_vec_15 = 1'b0;
    end
  end

  assign _zz_BTB_btb_write_index = (((((((BTB_btb_is_hit_vec_1 || BTB_btb_is_hit_vec_3) || BTB_btb_is_hit_vec_5) || BTB_btb_is_hit_vec_7) || BTB_btb_is_hit_vec_9) || BTB_btb_is_hit_vec_11) || BTB_btb_is_hit_vec_13) || BTB_btb_is_hit_vec_15);
  assign _zz_BTB_btb_write_index_1 = (((((((BTB_btb_is_hit_vec_2 || BTB_btb_is_hit_vec_3) || BTB_btb_is_hit_vec_6) || BTB_btb_is_hit_vec_7) || BTB_btb_is_hit_vec_10) || BTB_btb_is_hit_vec_11) || BTB_btb_is_hit_vec_14) || BTB_btb_is_hit_vec_15);
  assign _zz_BTB_btb_write_index_2 = (((((((BTB_btb_is_hit_vec_4 || BTB_btb_is_hit_vec_5) || BTB_btb_is_hit_vec_6) || BTB_btb_is_hit_vec_7) || BTB_btb_is_hit_vec_12) || BTB_btb_is_hit_vec_13) || BTB_btb_is_hit_vec_14) || BTB_btb_is_hit_vec_15);
  assign _zz_BTB_btb_write_index_3 = (((((((BTB_btb_is_hit_vec_8 || BTB_btb_is_hit_vec_9) || BTB_btb_is_hit_vec_10) || BTB_btb_is_hit_vec_11) || BTB_btb_is_hit_vec_12) || BTB_btb_is_hit_vec_13) || BTB_btb_is_hit_vec_14) || BTB_btb_is_hit_vec_15);
  assign BTB_btb_write_index = {_zz_BTB_btb_write_index_3,{_zz_BTB_btb_write_index_2,{_zz_BTB_btb_write_index_1,_zz_BTB_btb_write_index}}};
  assign _zz_34 = ({15'd0,1'b1} <<< BTB_btb_write_index);
  assign _zz_35 = ({15'd0,1'b1} <<< BTB_btb_write_index);
  assign _zz_36 = ({15'd0,1'b1} <<< BTB_btb_alloc_index_value);
  assign _zz_37 = ({15'd0,1'b1} <<< BTB_btb_alloc_index_value);
  assign RAS_ras_call_matched = (BTB_is_matched && BTB_is_call);
  assign RAS_ras_ret_matched = (BTB_is_matched && BTB_is_ret);
  assign when_Predictor_l169 = (train_valid && train_is_call);
  always @(*) begin
    if(when_Predictor_l169) begin
      RAS_ras_next_index_proven = (RAS_ras_curr_index_proven + 5'h01);
    end else begin
      if(when_Predictor_l172) begin
        RAS_ras_next_index_proven = (RAS_ras_curr_index_proven - 5'h01);
      end else begin
        RAS_ras_next_index_proven = RAS_ras_curr_index_proven;
      end
    end
  end

  assign when_Predictor_l172 = (train_valid && train_is_ret);
  assign when_Predictor_l180 = ((train_mispredicted && train_valid) && train_is_call);
  always @(*) begin
    if(when_Predictor_l180) begin
      RAS_ras_next_index = (RAS_ras_curr_index_proven + 5'h01);
    end else begin
      if(when_Predictor_l183) begin
        RAS_ras_next_index = (RAS_ras_curr_index_proven - 5'h01);
      end else begin
        if(RAS_ras_call_matched) begin
          RAS_ras_next_index = (RAS_ras_curr_index + 5'h01);
        end else begin
          if(RAS_ras_ret_matched) begin
            RAS_ras_next_index = (RAS_ras_curr_index - 5'h01);
          end else begin
            RAS_ras_next_index = RAS_ras_curr_index;
          end
        end
      end
    end
  end

  assign when_Predictor_l183 = ((train_mispredicted && train_valid) && train_is_ret);
  assign when_Predictor_l197 = ((train_mispredicted && train_valid) && train_is_call);
  assign _zz_38 = ({31'd0,1'b1} <<< RAS_ras_next_index);
  assign _zz_39 = _zz_38[0];
  assign _zz_40 = _zz_38[1];
  assign _zz_41 = _zz_38[2];
  assign _zz_42 = _zz_38[3];
  assign _zz_43 = _zz_38[4];
  assign _zz_44 = _zz_38[5];
  assign _zz_45 = _zz_38[6];
  assign _zz_46 = _zz_38[7];
  assign _zz_47 = _zz_38[8];
  assign _zz_48 = _zz_38[9];
  assign _zz_49 = _zz_38[10];
  assign _zz_50 = _zz_38[11];
  assign _zz_51 = _zz_38[12];
  assign _zz_52 = _zz_38[13];
  assign _zz_53 = _zz_38[14];
  assign _zz_54 = _zz_38[15];
  assign _zz_55 = _zz_38[16];
  assign _zz_56 = _zz_38[17];
  assign _zz_57 = _zz_38[18];
  assign _zz_58 = _zz_38[19];
  assign _zz_59 = _zz_38[20];
  assign _zz_60 = _zz_38[21];
  assign _zz_61 = _zz_38[22];
  assign _zz_62 = _zz_38[23];
  assign _zz_63 = _zz_38[24];
  assign _zz_64 = _zz_38[25];
  assign _zz_65 = _zz_38[26];
  assign _zz_66 = _zz_38[27];
  assign _zz_67 = _zz_38[28];
  assign _zz_68 = _zz_38[29];
  assign _zz_69 = _zz_38[30];
  assign _zz_70 = _zz_38[31];
  assign _zz_RAS_ras_regfile_0 = (train_pc + 64'h0000000000000004);
  assign _zz_RAS_ras_regfile_0_1 = (predict_pc + 64'h0000000000000004);
  assign when_Predictor_l205 = ((train_mispredicted && train_valid) && train_is_ret);
  assign RAS_ras_predict_pc = _zz_RAS_ras_predict_pc;
  assign predict_history = GSHARE_global_branch_history;
  assign predict_taken = (BTB_is_matched && (((GSHARE_pht_predict_taken || BTB_is_jmp) || BTB_is_call) || BTB_is_ret));
  assign predict_pc_next = (RAS_ras_ret_matched ? RAS_ras_predict_pc : ((BTB_is_matched && ((GSHARE_pht_predict_taken || BTB_is_jmp) || BTB_is_call)) ? BTB_target_pc_read : _zz_predict_pc_next));
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      GSHARE_global_branch_history <= 5'h0;
      GSHARE_PHT_0 <= 2'b01;
      GSHARE_PHT_1 <= 2'b01;
      GSHARE_PHT_2 <= 2'b01;
      GSHARE_PHT_3 <= 2'b01;
      GSHARE_PHT_4 <= 2'b01;
      GSHARE_PHT_5 <= 2'b01;
      GSHARE_PHT_6 <= 2'b01;
      GSHARE_PHT_7 <= 2'b01;
      GSHARE_PHT_8 <= 2'b01;
      GSHARE_PHT_9 <= 2'b01;
      GSHARE_PHT_10 <= 2'b01;
      GSHARE_PHT_11 <= 2'b01;
      GSHARE_PHT_12 <= 2'b01;
      GSHARE_PHT_13 <= 2'b01;
      GSHARE_PHT_14 <= 2'b01;
      GSHARE_PHT_15 <= 2'b01;
      GSHARE_PHT_16 <= 2'b01;
      GSHARE_PHT_17 <= 2'b01;
      GSHARE_PHT_18 <= 2'b01;
      GSHARE_PHT_19 <= 2'b01;
      GSHARE_PHT_20 <= 2'b01;
      GSHARE_PHT_21 <= 2'b01;
      GSHARE_PHT_22 <= 2'b01;
      GSHARE_PHT_23 <= 2'b01;
      GSHARE_PHT_24 <= 2'b01;
      GSHARE_PHT_25 <= 2'b01;
      GSHARE_PHT_26 <= 2'b01;
      GSHARE_PHT_27 <= 2'b01;
      GSHARE_PHT_28 <= 2'b01;
      GSHARE_PHT_29 <= 2'b01;
      GSHARE_PHT_30 <= 2'b01;
      GSHARE_PHT_31 <= 2'b01;
      BTB_valid <= 16'h0;
      BTB_source_pc_0 <= 64'h0;
      BTB_source_pc_1 <= 64'h0;
      BTB_source_pc_2 <= 64'h0;
      BTB_source_pc_3 <= 64'h0;
      BTB_source_pc_4 <= 64'h0;
      BTB_source_pc_5 <= 64'h0;
      BTB_source_pc_6 <= 64'h0;
      BTB_source_pc_7 <= 64'h0;
      BTB_source_pc_8 <= 64'h0;
      BTB_source_pc_9 <= 64'h0;
      BTB_source_pc_10 <= 64'h0;
      BTB_source_pc_11 <= 64'h0;
      BTB_source_pc_12 <= 64'h0;
      BTB_source_pc_13 <= 64'h0;
      BTB_source_pc_14 <= 64'h0;
      BTB_source_pc_15 <= 64'h0;
      BTB_call <= 16'h0;
      BTB_ret <= 16'h0;
      BTB_jmp <= 16'h0;
      BTB_target_pc_0 <= 64'h0;
      BTB_target_pc_1 <= 64'h0;
      BTB_target_pc_2 <= 64'h0;
      BTB_target_pc_3 <= 64'h0;
      BTB_target_pc_4 <= 64'h0;
      BTB_target_pc_5 <= 64'h0;
      BTB_target_pc_6 <= 64'h0;
      BTB_target_pc_7 <= 64'h0;
      BTB_target_pc_8 <= 64'h0;
      BTB_target_pc_9 <= 64'h0;
      BTB_target_pc_10 <= 64'h0;
      BTB_target_pc_11 <= 64'h0;
      BTB_target_pc_12 <= 64'h0;
      BTB_target_pc_13 <= 64'h0;
      BTB_target_pc_14 <= 64'h0;
      BTB_target_pc_15 <= 64'h0;
      BTB_btb_alloc_index_value <= 4'b0000;
      RAS_ras_curr_index <= 5'h0;
      RAS_ras_curr_index_proven <= 5'h0;
    end else begin
      if(train_valid) begin
        case(switch_Predictor_l38)
          2'b00 : begin
            if(train_taken) begin
              if(_zz_2) begin
                GSHARE_PHT_0 <= 2'b01;
              end
              if(_zz_3) begin
                GSHARE_PHT_1 <= 2'b01;
              end
              if(_zz_4) begin
                GSHARE_PHT_2 <= 2'b01;
              end
              if(_zz_5) begin
                GSHARE_PHT_3 <= 2'b01;
              end
              if(_zz_6) begin
                GSHARE_PHT_4 <= 2'b01;
              end
              if(_zz_7) begin
                GSHARE_PHT_5 <= 2'b01;
              end
              if(_zz_8) begin
                GSHARE_PHT_6 <= 2'b01;
              end
              if(_zz_9) begin
                GSHARE_PHT_7 <= 2'b01;
              end
              if(_zz_10) begin
                GSHARE_PHT_8 <= 2'b01;
              end
              if(_zz_11) begin
                GSHARE_PHT_9 <= 2'b01;
              end
              if(_zz_12) begin
                GSHARE_PHT_10 <= 2'b01;
              end
              if(_zz_13) begin
                GSHARE_PHT_11 <= 2'b01;
              end
              if(_zz_14) begin
                GSHARE_PHT_12 <= 2'b01;
              end
              if(_zz_15) begin
                GSHARE_PHT_13 <= 2'b01;
              end
              if(_zz_16) begin
                GSHARE_PHT_14 <= 2'b01;
              end
              if(_zz_17) begin
                GSHARE_PHT_15 <= 2'b01;
              end
              if(_zz_18) begin
                GSHARE_PHT_16 <= 2'b01;
              end
              if(_zz_19) begin
                GSHARE_PHT_17 <= 2'b01;
              end
              if(_zz_20) begin
                GSHARE_PHT_18 <= 2'b01;
              end
              if(_zz_21) begin
                GSHARE_PHT_19 <= 2'b01;
              end
              if(_zz_22) begin
                GSHARE_PHT_20 <= 2'b01;
              end
              if(_zz_23) begin
                GSHARE_PHT_21 <= 2'b01;
              end
              if(_zz_24) begin
                GSHARE_PHT_22 <= 2'b01;
              end
              if(_zz_25) begin
                GSHARE_PHT_23 <= 2'b01;
              end
              if(_zz_26) begin
                GSHARE_PHT_24 <= 2'b01;
              end
              if(_zz_27) begin
                GSHARE_PHT_25 <= 2'b01;
              end
              if(_zz_28) begin
                GSHARE_PHT_26 <= 2'b01;
              end
              if(_zz_29) begin
                GSHARE_PHT_27 <= 2'b01;
              end
              if(_zz_30) begin
                GSHARE_PHT_28 <= 2'b01;
              end
              if(_zz_31) begin
                GSHARE_PHT_29 <= 2'b01;
              end
              if(_zz_32) begin
                GSHARE_PHT_30 <= 2'b01;
              end
              if(_zz_33) begin
                GSHARE_PHT_31 <= 2'b01;
              end
            end else begin
              if(_zz_2) begin
                GSHARE_PHT_0 <= 2'b00;
              end
              if(_zz_3) begin
                GSHARE_PHT_1 <= 2'b00;
              end
              if(_zz_4) begin
                GSHARE_PHT_2 <= 2'b00;
              end
              if(_zz_5) begin
                GSHARE_PHT_3 <= 2'b00;
              end
              if(_zz_6) begin
                GSHARE_PHT_4 <= 2'b00;
              end
              if(_zz_7) begin
                GSHARE_PHT_5 <= 2'b00;
              end
              if(_zz_8) begin
                GSHARE_PHT_6 <= 2'b00;
              end
              if(_zz_9) begin
                GSHARE_PHT_7 <= 2'b00;
              end
              if(_zz_10) begin
                GSHARE_PHT_8 <= 2'b00;
              end
              if(_zz_11) begin
                GSHARE_PHT_9 <= 2'b00;
              end
              if(_zz_12) begin
                GSHARE_PHT_10 <= 2'b00;
              end
              if(_zz_13) begin
                GSHARE_PHT_11 <= 2'b00;
              end
              if(_zz_14) begin
                GSHARE_PHT_12 <= 2'b00;
              end
              if(_zz_15) begin
                GSHARE_PHT_13 <= 2'b00;
              end
              if(_zz_16) begin
                GSHARE_PHT_14 <= 2'b00;
              end
              if(_zz_17) begin
                GSHARE_PHT_15 <= 2'b00;
              end
              if(_zz_18) begin
                GSHARE_PHT_16 <= 2'b00;
              end
              if(_zz_19) begin
                GSHARE_PHT_17 <= 2'b00;
              end
              if(_zz_20) begin
                GSHARE_PHT_18 <= 2'b00;
              end
              if(_zz_21) begin
                GSHARE_PHT_19 <= 2'b00;
              end
              if(_zz_22) begin
                GSHARE_PHT_20 <= 2'b00;
              end
              if(_zz_23) begin
                GSHARE_PHT_21 <= 2'b00;
              end
              if(_zz_24) begin
                GSHARE_PHT_22 <= 2'b00;
              end
              if(_zz_25) begin
                GSHARE_PHT_23 <= 2'b00;
              end
              if(_zz_26) begin
                GSHARE_PHT_24 <= 2'b00;
              end
              if(_zz_27) begin
                GSHARE_PHT_25 <= 2'b00;
              end
              if(_zz_28) begin
                GSHARE_PHT_26 <= 2'b00;
              end
              if(_zz_29) begin
                GSHARE_PHT_27 <= 2'b00;
              end
              if(_zz_30) begin
                GSHARE_PHT_28 <= 2'b00;
              end
              if(_zz_31) begin
                GSHARE_PHT_29 <= 2'b00;
              end
              if(_zz_32) begin
                GSHARE_PHT_30 <= 2'b00;
              end
              if(_zz_33) begin
                GSHARE_PHT_31 <= 2'b00;
              end
            end
          end
          2'b01 : begin
            if(train_taken) begin
              if(_zz_2) begin
                GSHARE_PHT_0 <= 2'b10;
              end
              if(_zz_3) begin
                GSHARE_PHT_1 <= 2'b10;
              end
              if(_zz_4) begin
                GSHARE_PHT_2 <= 2'b10;
              end
              if(_zz_5) begin
                GSHARE_PHT_3 <= 2'b10;
              end
              if(_zz_6) begin
                GSHARE_PHT_4 <= 2'b10;
              end
              if(_zz_7) begin
                GSHARE_PHT_5 <= 2'b10;
              end
              if(_zz_8) begin
                GSHARE_PHT_6 <= 2'b10;
              end
              if(_zz_9) begin
                GSHARE_PHT_7 <= 2'b10;
              end
              if(_zz_10) begin
                GSHARE_PHT_8 <= 2'b10;
              end
              if(_zz_11) begin
                GSHARE_PHT_9 <= 2'b10;
              end
              if(_zz_12) begin
                GSHARE_PHT_10 <= 2'b10;
              end
              if(_zz_13) begin
                GSHARE_PHT_11 <= 2'b10;
              end
              if(_zz_14) begin
                GSHARE_PHT_12 <= 2'b10;
              end
              if(_zz_15) begin
                GSHARE_PHT_13 <= 2'b10;
              end
              if(_zz_16) begin
                GSHARE_PHT_14 <= 2'b10;
              end
              if(_zz_17) begin
                GSHARE_PHT_15 <= 2'b10;
              end
              if(_zz_18) begin
                GSHARE_PHT_16 <= 2'b10;
              end
              if(_zz_19) begin
                GSHARE_PHT_17 <= 2'b10;
              end
              if(_zz_20) begin
                GSHARE_PHT_18 <= 2'b10;
              end
              if(_zz_21) begin
                GSHARE_PHT_19 <= 2'b10;
              end
              if(_zz_22) begin
                GSHARE_PHT_20 <= 2'b10;
              end
              if(_zz_23) begin
                GSHARE_PHT_21 <= 2'b10;
              end
              if(_zz_24) begin
                GSHARE_PHT_22 <= 2'b10;
              end
              if(_zz_25) begin
                GSHARE_PHT_23 <= 2'b10;
              end
              if(_zz_26) begin
                GSHARE_PHT_24 <= 2'b10;
              end
              if(_zz_27) begin
                GSHARE_PHT_25 <= 2'b10;
              end
              if(_zz_28) begin
                GSHARE_PHT_26 <= 2'b10;
              end
              if(_zz_29) begin
                GSHARE_PHT_27 <= 2'b10;
              end
              if(_zz_30) begin
                GSHARE_PHT_28 <= 2'b10;
              end
              if(_zz_31) begin
                GSHARE_PHT_29 <= 2'b10;
              end
              if(_zz_32) begin
                GSHARE_PHT_30 <= 2'b10;
              end
              if(_zz_33) begin
                GSHARE_PHT_31 <= 2'b10;
              end
            end else begin
              if(_zz_2) begin
                GSHARE_PHT_0 <= 2'b00;
              end
              if(_zz_3) begin
                GSHARE_PHT_1 <= 2'b00;
              end
              if(_zz_4) begin
                GSHARE_PHT_2 <= 2'b00;
              end
              if(_zz_5) begin
                GSHARE_PHT_3 <= 2'b00;
              end
              if(_zz_6) begin
                GSHARE_PHT_4 <= 2'b00;
              end
              if(_zz_7) begin
                GSHARE_PHT_5 <= 2'b00;
              end
              if(_zz_8) begin
                GSHARE_PHT_6 <= 2'b00;
              end
              if(_zz_9) begin
                GSHARE_PHT_7 <= 2'b00;
              end
              if(_zz_10) begin
                GSHARE_PHT_8 <= 2'b00;
              end
              if(_zz_11) begin
                GSHARE_PHT_9 <= 2'b00;
              end
              if(_zz_12) begin
                GSHARE_PHT_10 <= 2'b00;
              end
              if(_zz_13) begin
                GSHARE_PHT_11 <= 2'b00;
              end
              if(_zz_14) begin
                GSHARE_PHT_12 <= 2'b00;
              end
              if(_zz_15) begin
                GSHARE_PHT_13 <= 2'b00;
              end
              if(_zz_16) begin
                GSHARE_PHT_14 <= 2'b00;
              end
              if(_zz_17) begin
                GSHARE_PHT_15 <= 2'b00;
              end
              if(_zz_18) begin
                GSHARE_PHT_16 <= 2'b00;
              end
              if(_zz_19) begin
                GSHARE_PHT_17 <= 2'b00;
              end
              if(_zz_20) begin
                GSHARE_PHT_18 <= 2'b00;
              end
              if(_zz_21) begin
                GSHARE_PHT_19 <= 2'b00;
              end
              if(_zz_22) begin
                GSHARE_PHT_20 <= 2'b00;
              end
              if(_zz_23) begin
                GSHARE_PHT_21 <= 2'b00;
              end
              if(_zz_24) begin
                GSHARE_PHT_22 <= 2'b00;
              end
              if(_zz_25) begin
                GSHARE_PHT_23 <= 2'b00;
              end
              if(_zz_26) begin
                GSHARE_PHT_24 <= 2'b00;
              end
              if(_zz_27) begin
                GSHARE_PHT_25 <= 2'b00;
              end
              if(_zz_28) begin
                GSHARE_PHT_26 <= 2'b00;
              end
              if(_zz_29) begin
                GSHARE_PHT_27 <= 2'b00;
              end
              if(_zz_30) begin
                GSHARE_PHT_28 <= 2'b00;
              end
              if(_zz_31) begin
                GSHARE_PHT_29 <= 2'b00;
              end
              if(_zz_32) begin
                GSHARE_PHT_30 <= 2'b00;
              end
              if(_zz_33) begin
                GSHARE_PHT_31 <= 2'b00;
              end
            end
          end
          2'b10 : begin
            if(train_taken) begin
              if(_zz_2) begin
                GSHARE_PHT_0 <= 2'b11;
              end
              if(_zz_3) begin
                GSHARE_PHT_1 <= 2'b11;
              end
              if(_zz_4) begin
                GSHARE_PHT_2 <= 2'b11;
              end
              if(_zz_5) begin
                GSHARE_PHT_3 <= 2'b11;
              end
              if(_zz_6) begin
                GSHARE_PHT_4 <= 2'b11;
              end
              if(_zz_7) begin
                GSHARE_PHT_5 <= 2'b11;
              end
              if(_zz_8) begin
                GSHARE_PHT_6 <= 2'b11;
              end
              if(_zz_9) begin
                GSHARE_PHT_7 <= 2'b11;
              end
              if(_zz_10) begin
                GSHARE_PHT_8 <= 2'b11;
              end
              if(_zz_11) begin
                GSHARE_PHT_9 <= 2'b11;
              end
              if(_zz_12) begin
                GSHARE_PHT_10 <= 2'b11;
              end
              if(_zz_13) begin
                GSHARE_PHT_11 <= 2'b11;
              end
              if(_zz_14) begin
                GSHARE_PHT_12 <= 2'b11;
              end
              if(_zz_15) begin
                GSHARE_PHT_13 <= 2'b11;
              end
              if(_zz_16) begin
                GSHARE_PHT_14 <= 2'b11;
              end
              if(_zz_17) begin
                GSHARE_PHT_15 <= 2'b11;
              end
              if(_zz_18) begin
                GSHARE_PHT_16 <= 2'b11;
              end
              if(_zz_19) begin
                GSHARE_PHT_17 <= 2'b11;
              end
              if(_zz_20) begin
                GSHARE_PHT_18 <= 2'b11;
              end
              if(_zz_21) begin
                GSHARE_PHT_19 <= 2'b11;
              end
              if(_zz_22) begin
                GSHARE_PHT_20 <= 2'b11;
              end
              if(_zz_23) begin
                GSHARE_PHT_21 <= 2'b11;
              end
              if(_zz_24) begin
                GSHARE_PHT_22 <= 2'b11;
              end
              if(_zz_25) begin
                GSHARE_PHT_23 <= 2'b11;
              end
              if(_zz_26) begin
                GSHARE_PHT_24 <= 2'b11;
              end
              if(_zz_27) begin
                GSHARE_PHT_25 <= 2'b11;
              end
              if(_zz_28) begin
                GSHARE_PHT_26 <= 2'b11;
              end
              if(_zz_29) begin
                GSHARE_PHT_27 <= 2'b11;
              end
              if(_zz_30) begin
                GSHARE_PHT_28 <= 2'b11;
              end
              if(_zz_31) begin
                GSHARE_PHT_29 <= 2'b11;
              end
              if(_zz_32) begin
                GSHARE_PHT_30 <= 2'b11;
              end
              if(_zz_33) begin
                GSHARE_PHT_31 <= 2'b11;
              end
            end else begin
              if(_zz_2) begin
                GSHARE_PHT_0 <= 2'b00;
              end
              if(_zz_3) begin
                GSHARE_PHT_1 <= 2'b00;
              end
              if(_zz_4) begin
                GSHARE_PHT_2 <= 2'b00;
              end
              if(_zz_5) begin
                GSHARE_PHT_3 <= 2'b00;
              end
              if(_zz_6) begin
                GSHARE_PHT_4 <= 2'b00;
              end
              if(_zz_7) begin
                GSHARE_PHT_5 <= 2'b00;
              end
              if(_zz_8) begin
                GSHARE_PHT_6 <= 2'b00;
              end
              if(_zz_9) begin
                GSHARE_PHT_7 <= 2'b00;
              end
              if(_zz_10) begin
                GSHARE_PHT_8 <= 2'b00;
              end
              if(_zz_11) begin
                GSHARE_PHT_9 <= 2'b00;
              end
              if(_zz_12) begin
                GSHARE_PHT_10 <= 2'b00;
              end
              if(_zz_13) begin
                GSHARE_PHT_11 <= 2'b00;
              end
              if(_zz_14) begin
                GSHARE_PHT_12 <= 2'b00;
              end
              if(_zz_15) begin
                GSHARE_PHT_13 <= 2'b00;
              end
              if(_zz_16) begin
                GSHARE_PHT_14 <= 2'b00;
              end
              if(_zz_17) begin
                GSHARE_PHT_15 <= 2'b00;
              end
              if(_zz_18) begin
                GSHARE_PHT_16 <= 2'b00;
              end
              if(_zz_19) begin
                GSHARE_PHT_17 <= 2'b00;
              end
              if(_zz_20) begin
                GSHARE_PHT_18 <= 2'b00;
              end
              if(_zz_21) begin
                GSHARE_PHT_19 <= 2'b00;
              end
              if(_zz_22) begin
                GSHARE_PHT_20 <= 2'b00;
              end
              if(_zz_23) begin
                GSHARE_PHT_21 <= 2'b00;
              end
              if(_zz_24) begin
                GSHARE_PHT_22 <= 2'b00;
              end
              if(_zz_25) begin
                GSHARE_PHT_23 <= 2'b00;
              end
              if(_zz_26) begin
                GSHARE_PHT_24 <= 2'b00;
              end
              if(_zz_27) begin
                GSHARE_PHT_25 <= 2'b00;
              end
              if(_zz_28) begin
                GSHARE_PHT_26 <= 2'b00;
              end
              if(_zz_29) begin
                GSHARE_PHT_27 <= 2'b00;
              end
              if(_zz_30) begin
                GSHARE_PHT_28 <= 2'b00;
              end
              if(_zz_31) begin
                GSHARE_PHT_29 <= 2'b00;
              end
              if(_zz_32) begin
                GSHARE_PHT_30 <= 2'b00;
              end
              if(_zz_33) begin
                GSHARE_PHT_31 <= 2'b00;
              end
            end
          end
          default : begin
            if(when_Predictor_l61) begin
              if(_zz_2) begin
                GSHARE_PHT_0 <= 2'b10;
              end
              if(_zz_3) begin
                GSHARE_PHT_1 <= 2'b10;
              end
              if(_zz_4) begin
                GSHARE_PHT_2 <= 2'b10;
              end
              if(_zz_5) begin
                GSHARE_PHT_3 <= 2'b10;
              end
              if(_zz_6) begin
                GSHARE_PHT_4 <= 2'b10;
              end
              if(_zz_7) begin
                GSHARE_PHT_5 <= 2'b10;
              end
              if(_zz_8) begin
                GSHARE_PHT_6 <= 2'b10;
              end
              if(_zz_9) begin
                GSHARE_PHT_7 <= 2'b10;
              end
              if(_zz_10) begin
                GSHARE_PHT_8 <= 2'b10;
              end
              if(_zz_11) begin
                GSHARE_PHT_9 <= 2'b10;
              end
              if(_zz_12) begin
                GSHARE_PHT_10 <= 2'b10;
              end
              if(_zz_13) begin
                GSHARE_PHT_11 <= 2'b10;
              end
              if(_zz_14) begin
                GSHARE_PHT_12 <= 2'b10;
              end
              if(_zz_15) begin
                GSHARE_PHT_13 <= 2'b10;
              end
              if(_zz_16) begin
                GSHARE_PHT_14 <= 2'b10;
              end
              if(_zz_17) begin
                GSHARE_PHT_15 <= 2'b10;
              end
              if(_zz_18) begin
                GSHARE_PHT_16 <= 2'b10;
              end
              if(_zz_19) begin
                GSHARE_PHT_17 <= 2'b10;
              end
              if(_zz_20) begin
                GSHARE_PHT_18 <= 2'b10;
              end
              if(_zz_21) begin
                GSHARE_PHT_19 <= 2'b10;
              end
              if(_zz_22) begin
                GSHARE_PHT_20 <= 2'b10;
              end
              if(_zz_23) begin
                GSHARE_PHT_21 <= 2'b10;
              end
              if(_zz_24) begin
                GSHARE_PHT_22 <= 2'b10;
              end
              if(_zz_25) begin
                GSHARE_PHT_23 <= 2'b10;
              end
              if(_zz_26) begin
                GSHARE_PHT_24 <= 2'b10;
              end
              if(_zz_27) begin
                GSHARE_PHT_25 <= 2'b10;
              end
              if(_zz_28) begin
                GSHARE_PHT_26 <= 2'b10;
              end
              if(_zz_29) begin
                GSHARE_PHT_27 <= 2'b10;
              end
              if(_zz_30) begin
                GSHARE_PHT_28 <= 2'b10;
              end
              if(_zz_31) begin
                GSHARE_PHT_29 <= 2'b10;
              end
              if(_zz_32) begin
                GSHARE_PHT_30 <= 2'b10;
              end
              if(_zz_33) begin
                GSHARE_PHT_31 <= 2'b10;
              end
            end else begin
              if(_zz_2) begin
                GSHARE_PHT_0 <= 2'b11;
              end
              if(_zz_3) begin
                GSHARE_PHT_1 <= 2'b11;
              end
              if(_zz_4) begin
                GSHARE_PHT_2 <= 2'b11;
              end
              if(_zz_5) begin
                GSHARE_PHT_3 <= 2'b11;
              end
              if(_zz_6) begin
                GSHARE_PHT_4 <= 2'b11;
              end
              if(_zz_7) begin
                GSHARE_PHT_5 <= 2'b11;
              end
              if(_zz_8) begin
                GSHARE_PHT_6 <= 2'b11;
              end
              if(_zz_9) begin
                GSHARE_PHT_7 <= 2'b11;
              end
              if(_zz_10) begin
                GSHARE_PHT_8 <= 2'b11;
              end
              if(_zz_11) begin
                GSHARE_PHT_9 <= 2'b11;
              end
              if(_zz_12) begin
                GSHARE_PHT_10 <= 2'b11;
              end
              if(_zz_13) begin
                GSHARE_PHT_11 <= 2'b11;
              end
              if(_zz_14) begin
                GSHARE_PHT_12 <= 2'b11;
              end
              if(_zz_15) begin
                GSHARE_PHT_13 <= 2'b11;
              end
              if(_zz_16) begin
                GSHARE_PHT_14 <= 2'b11;
              end
              if(_zz_17) begin
                GSHARE_PHT_15 <= 2'b11;
              end
              if(_zz_18) begin
                GSHARE_PHT_16 <= 2'b11;
              end
              if(_zz_19) begin
                GSHARE_PHT_17 <= 2'b11;
              end
              if(_zz_20) begin
                GSHARE_PHT_18 <= 2'b11;
              end
              if(_zz_21) begin
                GSHARE_PHT_19 <= 2'b11;
              end
              if(_zz_22) begin
                GSHARE_PHT_20 <= 2'b11;
              end
              if(_zz_23) begin
                GSHARE_PHT_21 <= 2'b11;
              end
              if(_zz_24) begin
                GSHARE_PHT_22 <= 2'b11;
              end
              if(_zz_25) begin
                GSHARE_PHT_23 <= 2'b11;
              end
              if(_zz_26) begin
                GSHARE_PHT_24 <= 2'b11;
              end
              if(_zz_27) begin
                GSHARE_PHT_25 <= 2'b11;
              end
              if(_zz_28) begin
                GSHARE_PHT_26 <= 2'b11;
              end
              if(_zz_29) begin
                GSHARE_PHT_27 <= 2'b11;
              end
              if(_zz_30) begin
                GSHARE_PHT_28 <= 2'b11;
              end
              if(_zz_31) begin
                GSHARE_PHT_29 <= 2'b11;
              end
              if(_zz_32) begin
                GSHARE_PHT_30 <= 2'b11;
              end
              if(_zz_33) begin
                GSHARE_PHT_31 <= 2'b11;
              end
            end
          end
        endcase
      end
      if(when_Predictor_l70) begin
        GSHARE_global_branch_history <= {train_history[3 : 0],train_taken};
      end else begin
        if(predict_valid) begin
          GSHARE_global_branch_history <= {GSHARE_global_branch_history[3 : 0],predict_taken};
        end
      end
      BTB_btb_alloc_index_value <= BTB_btb_alloc_index_valueNext;
      if(BTB_btb_is_hit) begin
        if(_zz_34[0]) begin
          BTB_source_pc_0 <= train_pc;
        end
        if(_zz_34[1]) begin
          BTB_source_pc_1 <= train_pc;
        end
        if(_zz_34[2]) begin
          BTB_source_pc_2 <= train_pc;
        end
        if(_zz_34[3]) begin
          BTB_source_pc_3 <= train_pc;
        end
        if(_zz_34[4]) begin
          BTB_source_pc_4 <= train_pc;
        end
        if(_zz_34[5]) begin
          BTB_source_pc_5 <= train_pc;
        end
        if(_zz_34[6]) begin
          BTB_source_pc_6 <= train_pc;
        end
        if(_zz_34[7]) begin
          BTB_source_pc_7 <= train_pc;
        end
        if(_zz_34[8]) begin
          BTB_source_pc_8 <= train_pc;
        end
        if(_zz_34[9]) begin
          BTB_source_pc_9 <= train_pc;
        end
        if(_zz_34[10]) begin
          BTB_source_pc_10 <= train_pc;
        end
        if(_zz_34[11]) begin
          BTB_source_pc_11 <= train_pc;
        end
        if(_zz_34[12]) begin
          BTB_source_pc_12 <= train_pc;
        end
        if(_zz_34[13]) begin
          BTB_source_pc_13 <= train_pc;
        end
        if(_zz_34[14]) begin
          BTB_source_pc_14 <= train_pc;
        end
        if(_zz_34[15]) begin
          BTB_source_pc_15 <= train_pc;
        end
        BTB_call[BTB_btb_write_index] <= train_is_call;
        BTB_ret[BTB_btb_write_index] <= train_is_ret;
        BTB_jmp[BTB_btb_write_index] <= train_is_jmp;
        if(_zz_35[0]) begin
          BTB_target_pc_0 <= train_pc_next;
        end
        if(_zz_35[1]) begin
          BTB_target_pc_1 <= train_pc_next;
        end
        if(_zz_35[2]) begin
          BTB_target_pc_2 <= train_pc_next;
        end
        if(_zz_35[3]) begin
          BTB_target_pc_3 <= train_pc_next;
        end
        if(_zz_35[4]) begin
          BTB_target_pc_4 <= train_pc_next;
        end
        if(_zz_35[5]) begin
          BTB_target_pc_5 <= train_pc_next;
        end
        if(_zz_35[6]) begin
          BTB_target_pc_6 <= train_pc_next;
        end
        if(_zz_35[7]) begin
          BTB_target_pc_7 <= train_pc_next;
        end
        if(_zz_35[8]) begin
          BTB_target_pc_8 <= train_pc_next;
        end
        if(_zz_35[9]) begin
          BTB_target_pc_9 <= train_pc_next;
        end
        if(_zz_35[10]) begin
          BTB_target_pc_10 <= train_pc_next;
        end
        if(_zz_35[11]) begin
          BTB_target_pc_11 <= train_pc_next;
        end
        if(_zz_35[12]) begin
          BTB_target_pc_12 <= train_pc_next;
        end
        if(_zz_35[13]) begin
          BTB_target_pc_13 <= train_pc_next;
        end
        if(_zz_35[14]) begin
          BTB_target_pc_14 <= train_pc_next;
        end
        if(_zz_35[15]) begin
          BTB_target_pc_15 <= train_pc_next;
        end
      end else begin
        if(BTB_btb_is_miss) begin
          BTB_valid[BTB_btb_alloc_index_value] <= 1'b1;
          if(_zz_36[0]) begin
            BTB_source_pc_0 <= train_pc;
          end
          if(_zz_36[1]) begin
            BTB_source_pc_1 <= train_pc;
          end
          if(_zz_36[2]) begin
            BTB_source_pc_2 <= train_pc;
          end
          if(_zz_36[3]) begin
            BTB_source_pc_3 <= train_pc;
          end
          if(_zz_36[4]) begin
            BTB_source_pc_4 <= train_pc;
          end
          if(_zz_36[5]) begin
            BTB_source_pc_5 <= train_pc;
          end
          if(_zz_36[6]) begin
            BTB_source_pc_6 <= train_pc;
          end
          if(_zz_36[7]) begin
            BTB_source_pc_7 <= train_pc;
          end
          if(_zz_36[8]) begin
            BTB_source_pc_8 <= train_pc;
          end
          if(_zz_36[9]) begin
            BTB_source_pc_9 <= train_pc;
          end
          if(_zz_36[10]) begin
            BTB_source_pc_10 <= train_pc;
          end
          if(_zz_36[11]) begin
            BTB_source_pc_11 <= train_pc;
          end
          if(_zz_36[12]) begin
            BTB_source_pc_12 <= train_pc;
          end
          if(_zz_36[13]) begin
            BTB_source_pc_13 <= train_pc;
          end
          if(_zz_36[14]) begin
            BTB_source_pc_14 <= train_pc;
          end
          if(_zz_36[15]) begin
            BTB_source_pc_15 <= train_pc;
          end
          BTB_call[BTB_btb_alloc_index_value] <= train_is_call;
          BTB_ret[BTB_btb_alloc_index_value] <= train_is_ret;
          BTB_jmp[BTB_btb_alloc_index_value] <= train_is_jmp;
          if(_zz_37[0]) begin
            BTB_target_pc_0 <= train_pc_next;
          end
          if(_zz_37[1]) begin
            BTB_target_pc_1 <= train_pc_next;
          end
          if(_zz_37[2]) begin
            BTB_target_pc_2 <= train_pc_next;
          end
          if(_zz_37[3]) begin
            BTB_target_pc_3 <= train_pc_next;
          end
          if(_zz_37[4]) begin
            BTB_target_pc_4 <= train_pc_next;
          end
          if(_zz_37[5]) begin
            BTB_target_pc_5 <= train_pc_next;
          end
          if(_zz_37[6]) begin
            BTB_target_pc_6 <= train_pc_next;
          end
          if(_zz_37[7]) begin
            BTB_target_pc_7 <= train_pc_next;
          end
          if(_zz_37[8]) begin
            BTB_target_pc_8 <= train_pc_next;
          end
          if(_zz_37[9]) begin
            BTB_target_pc_9 <= train_pc_next;
          end
          if(_zz_37[10]) begin
            BTB_target_pc_10 <= train_pc_next;
          end
          if(_zz_37[11]) begin
            BTB_target_pc_11 <= train_pc_next;
          end
          if(_zz_37[12]) begin
            BTB_target_pc_12 <= train_pc_next;
          end
          if(_zz_37[13]) begin
            BTB_target_pc_13 <= train_pc_next;
          end
          if(_zz_37[14]) begin
            BTB_target_pc_14 <= train_pc_next;
          end
          if(_zz_37[15]) begin
            BTB_target_pc_15 <= train_pc_next;
          end
        end
      end
      RAS_ras_curr_index_proven <= RAS_ras_next_index;
      if(when_Predictor_l197) begin
        RAS_ras_curr_index <= RAS_ras_next_index;
      end else begin
        if(RAS_ras_call_matched) begin
          RAS_ras_curr_index <= RAS_ras_next_index;
        end else begin
          if(when_Predictor_l205) begin
            RAS_ras_curr_index <= RAS_ras_next_index;
          end else begin
            if(RAS_ras_ret_matched) begin
              RAS_ras_curr_index <= RAS_ras_next_index;
            end
          end
        end
      end
    end
  end

  always @(posedge io_axiClk) begin
    if(when_Predictor_l197) begin
      if(_zz_39) begin
        RAS_ras_regfile_0 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_40) begin
        RAS_ras_regfile_1 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_41) begin
        RAS_ras_regfile_2 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_42) begin
        RAS_ras_regfile_3 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_43) begin
        RAS_ras_regfile_4 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_44) begin
        RAS_ras_regfile_5 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_45) begin
        RAS_ras_regfile_6 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_46) begin
        RAS_ras_regfile_7 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_47) begin
        RAS_ras_regfile_8 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_48) begin
        RAS_ras_regfile_9 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_49) begin
        RAS_ras_regfile_10 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_50) begin
        RAS_ras_regfile_11 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_51) begin
        RAS_ras_regfile_12 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_52) begin
        RAS_ras_regfile_13 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_53) begin
        RAS_ras_regfile_14 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_54) begin
        RAS_ras_regfile_15 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_55) begin
        RAS_ras_regfile_16 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_56) begin
        RAS_ras_regfile_17 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_57) begin
        RAS_ras_regfile_18 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_58) begin
        RAS_ras_regfile_19 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_59) begin
        RAS_ras_regfile_20 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_60) begin
        RAS_ras_regfile_21 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_61) begin
        RAS_ras_regfile_22 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_62) begin
        RAS_ras_regfile_23 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_63) begin
        RAS_ras_regfile_24 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_64) begin
        RAS_ras_regfile_25 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_65) begin
        RAS_ras_regfile_26 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_66) begin
        RAS_ras_regfile_27 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_67) begin
        RAS_ras_regfile_28 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_68) begin
        RAS_ras_regfile_29 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_69) begin
        RAS_ras_regfile_30 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_70) begin
        RAS_ras_regfile_31 <= _zz_RAS_ras_regfile_0;
      end
    end else begin
      if(RAS_ras_call_matched) begin
        if(_zz_39) begin
          RAS_ras_regfile_0 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_40) begin
          RAS_ras_regfile_1 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_41) begin
          RAS_ras_regfile_2 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_42) begin
          RAS_ras_regfile_3 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_43) begin
          RAS_ras_regfile_4 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_44) begin
          RAS_ras_regfile_5 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_45) begin
          RAS_ras_regfile_6 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_46) begin
          RAS_ras_regfile_7 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_47) begin
          RAS_ras_regfile_8 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_48) begin
          RAS_ras_regfile_9 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_49) begin
          RAS_ras_regfile_10 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_50) begin
          RAS_ras_regfile_11 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_51) begin
          RAS_ras_regfile_12 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_52) begin
          RAS_ras_regfile_13 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_53) begin
          RAS_ras_regfile_14 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_54) begin
          RAS_ras_regfile_15 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_55) begin
          RAS_ras_regfile_16 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_56) begin
          RAS_ras_regfile_17 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_57) begin
          RAS_ras_regfile_18 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_58) begin
          RAS_ras_regfile_19 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_59) begin
          RAS_ras_regfile_20 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_60) begin
          RAS_ras_regfile_21 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_61) begin
          RAS_ras_regfile_22 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_62) begin
          RAS_ras_regfile_23 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_63) begin
          RAS_ras_regfile_24 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_64) begin
          RAS_ras_regfile_25 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_65) begin
          RAS_ras_regfile_26 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_66) begin
          RAS_ras_regfile_27 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_67) begin
          RAS_ras_regfile_28 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_68) begin
          RAS_ras_regfile_29 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_69) begin
          RAS_ras_regfile_30 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_70) begin
          RAS_ras_regfile_31 <= _zz_RAS_ras_regfile_0_1;
        end
      end
    end
  end


endmodule

module FIFO_2 (
  input               ports_s_ports_valid,
  output              ports_s_ports_ready,
  input      [31:0]   ports_s_ports_payload,
  output              ports_m_ports_valid,
  input               ports_m_ports_ready,
  output     [31:0]   ports_m_ports_payload,
  input               flush,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  reg        [31:0]   _zz_ports_m_ports_payload;
  reg        [2:0]    read_ptr;
  reg        [2:0]    write_ptr;
  wire       [1:0]    read_addr;
  wire       [1:0]    next_read_addr;
  wire       [1:0]    write_addr;
  wire                fifo_empty;
  wire                fifo_full;
  reg        [31:0]   fifo_ram_0;
  reg        [31:0]   fifo_ram_1;
  reg        [31:0]   fifo_ram_2;
  reg        [31:0]   fifo_ram_3;
  wire                ports_m_ports_fire;
  wire       [3:0]    _zz_1;
  wire                ports_s_ports_fire;

  always @(*) begin
    case(read_addr)
      2'b00 : _zz_ports_m_ports_payload = fifo_ram_0;
      2'b01 : _zz_ports_m_ports_payload = fifo_ram_1;
      2'b10 : _zz_ports_m_ports_payload = fifo_ram_2;
      default : _zz_ports_m_ports_payload = fifo_ram_3;
    endcase
  end

  assign read_addr = read_ptr[1 : 0];
  assign next_read_addr = (read_addr + 2'b01);
  assign write_addr = write_ptr[1 : 0];
  assign fifo_empty = (read_ptr == write_ptr);
  assign fifo_full = ((read_addr == write_addr) && (read_ptr[2] != write_ptr[2]));
  assign ports_m_ports_fire = (ports_m_ports_valid && ports_m_ports_ready);
  assign _zz_1 = ({3'd0,1'b1} <<< write_addr);
  assign ports_s_ports_fire = (ports_s_ports_valid && ports_s_ports_ready);
  assign ports_s_ports_ready = (! fifo_full);
  assign ports_m_ports_valid = (! fifo_empty);
  assign ports_m_ports_payload = _zz_ports_m_ports_payload;
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      read_ptr <= 3'b000;
      write_ptr <= 3'b000;
    end else begin
      if(flush) begin
        read_ptr <= 3'b000;
      end else begin
        if(ports_m_ports_fire) begin
          read_ptr <= (read_ptr + 3'b001);
        end
      end
      if(flush) begin
        write_ptr <= 3'b000;
      end else begin
        if(ports_s_ports_fire) begin
          write_ptr <= (write_ptr + 3'b001);
        end
      end
    end
  end

  always @(posedge io_axiClk) begin
    if(!flush) begin
      if(ports_s_ports_fire) begin
        if(_zz_1[0]) begin
          fifo_ram_0 <= ports_s_ports_payload;
        end
        if(_zz_1[1]) begin
          fifo_ram_1 <= ports_s_ports_payload;
        end
        if(_zz_1[2]) begin
          fifo_ram_2 <= ports_s_ports_payload;
        end
        if(_zz_1[3]) begin
          fifo_ram_3 <= ports_s_ports_payload;
        end
      end
    end
  end


endmodule

module FIFO_1 (
  input               ports_s_ports_valid,
  output              ports_s_ports_ready,
  input               ports_s_ports_payload,
  output              ports_m_ports_valid,
  input               ports_m_ports_ready,
  output              ports_m_ports_payload,
  input               flush,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  reg                 _zz_ports_m_ports_payload;
  reg        [2:0]    read_ptr;
  reg        [2:0]    write_ptr;
  wire       [1:0]    read_addr;
  wire       [1:0]    next_read_addr;
  wire       [1:0]    write_addr;
  wire                fifo_empty;
  wire                fifo_full;
  reg                 fifo_ram_0;
  reg                 fifo_ram_1;
  reg                 fifo_ram_2;
  reg                 fifo_ram_3;
  wire                ports_m_ports_fire;
  wire       [3:0]    _zz_1;
  wire                ports_s_ports_fire;

  always @(*) begin
    case(read_addr)
      2'b00 : _zz_ports_m_ports_payload = fifo_ram_0;
      2'b01 : _zz_ports_m_ports_payload = fifo_ram_1;
      2'b10 : _zz_ports_m_ports_payload = fifo_ram_2;
      default : _zz_ports_m_ports_payload = fifo_ram_3;
    endcase
  end

  assign read_addr = read_ptr[1 : 0];
  assign next_read_addr = (read_addr + 2'b01);
  assign write_addr = write_ptr[1 : 0];
  assign fifo_empty = (read_ptr == write_ptr);
  assign fifo_full = ((read_addr == write_addr) && (read_ptr[2] != write_ptr[2]));
  assign ports_m_ports_fire = (ports_m_ports_valid && ports_m_ports_ready);
  assign _zz_1 = ({3'd0,1'b1} <<< write_addr);
  assign ports_s_ports_fire = (ports_s_ports_valid && ports_s_ports_ready);
  assign ports_s_ports_ready = (! fifo_full);
  assign ports_m_ports_valid = (! fifo_empty);
  assign ports_m_ports_payload = _zz_ports_m_ports_payload;
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      read_ptr <= 3'b000;
      write_ptr <= 3'b000;
    end else begin
      if(flush) begin
        read_ptr <= 3'b000;
      end else begin
        if(ports_m_ports_fire) begin
          read_ptr <= (read_ptr + 3'b001);
        end
      end
      if(flush) begin
        write_ptr <= 3'b000;
      end else begin
        if(ports_s_ports_fire) begin
          write_ptr <= (write_ptr + 3'b001);
        end
      end
    end
  end

  always @(posedge io_axiClk) begin
    if(!flush) begin
      if(ports_s_ports_fire) begin
        if(_zz_1[0]) begin
          fifo_ram_0 <= ports_s_ports_payload;
        end
        if(_zz_1[1]) begin
          fifo_ram_1 <= ports_s_ports_payload;
        end
        if(_zz_1[2]) begin
          fifo_ram_2 <= ports_s_ports_payload;
        end
        if(_zz_1[3]) begin
          fifo_ram_3 <= ports_s_ports_payload;
        end
      end
    end
  end


endmodule

module FIFO (
  input               ports_s_ports_valid,
  output              ports_s_ports_ready,
  input      [63:0]   ports_s_ports_payload,
  output              ports_m_ports_valid,
  input               ports_m_ports_ready,
  output     [63:0]   ports_m_ports_payload,
  input               flush,
  output     [63:0]   next_payload,
  output              next_valid,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  reg        [63:0]   _zz_ports_m_ports_payload;
  reg        [63:0]   _zz_next_payload;
  reg        [2:0]    read_ptr;
  reg        [2:0]    write_ptr;
  wire       [1:0]    read_addr;
  wire       [1:0]    next_read_addr;
  wire       [1:0]    write_addr;
  wire                fifo_empty;
  wire                fifo_full;
  reg        [63:0]   fifo_ram_0;
  reg        [63:0]   fifo_ram_1;
  reg        [63:0]   fifo_ram_2;
  reg        [63:0]   fifo_ram_3;
  wire                ports_m_ports_fire;
  wire       [3:0]    _zz_1;
  wire                ports_s_ports_fire;
  reg        [2:0]    fifo_cnt;
  wire                ports_s_ports_fire_1;
  wire                ports_m_ports_fire_1;
  wire                when_FIFO_l61;
  wire                ports_s_ports_fire_2;
  wire                ports_m_ports_fire_2;
  wire                when_FIFO_l64;

  always @(*) begin
    case(read_addr)
      2'b00 : _zz_ports_m_ports_payload = fifo_ram_0;
      2'b01 : _zz_ports_m_ports_payload = fifo_ram_1;
      2'b10 : _zz_ports_m_ports_payload = fifo_ram_2;
      default : _zz_ports_m_ports_payload = fifo_ram_3;
    endcase
  end

  always @(*) begin
    case(next_read_addr)
      2'b00 : _zz_next_payload = fifo_ram_0;
      2'b01 : _zz_next_payload = fifo_ram_1;
      2'b10 : _zz_next_payload = fifo_ram_2;
      default : _zz_next_payload = fifo_ram_3;
    endcase
  end

  assign read_addr = read_ptr[1 : 0];
  assign next_read_addr = (read_addr + 2'b01);
  assign write_addr = write_ptr[1 : 0];
  assign fifo_empty = (read_ptr == write_ptr);
  assign fifo_full = ((read_addr == write_addr) && (read_ptr[2] != write_ptr[2]));
  assign ports_m_ports_fire = (ports_m_ports_valid && ports_m_ports_ready);
  assign _zz_1 = ({3'd0,1'b1} <<< write_addr);
  assign ports_s_ports_fire = (ports_s_ports_valid && ports_s_ports_ready);
  assign ports_s_ports_ready = (! fifo_full);
  assign ports_m_ports_valid = (! fifo_empty);
  assign ports_m_ports_payload = _zz_ports_m_ports_payload;
  assign next_payload = _zz_next_payload;
  assign ports_s_ports_fire_1 = (ports_s_ports_valid && ports_s_ports_ready);
  assign ports_m_ports_fire_1 = (ports_m_ports_valid && ports_m_ports_ready);
  assign when_FIFO_l61 = (ports_s_ports_fire_1 && (! ports_m_ports_fire_1));
  assign ports_s_ports_fire_2 = (ports_s_ports_valid && ports_s_ports_ready);
  assign ports_m_ports_fire_2 = (ports_m_ports_valid && ports_m_ports_ready);
  assign when_FIFO_l64 = ((! ports_s_ports_fire_2) && ports_m_ports_fire_2);
  assign next_valid = (3'b010 <= fifo_cnt);
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      read_ptr <= 3'b000;
      write_ptr <= 3'b000;
      fifo_cnt <= 3'b000;
    end else begin
      if(flush) begin
        read_ptr <= 3'b000;
      end else begin
        if(ports_m_ports_fire) begin
          read_ptr <= (read_ptr + 3'b001);
        end
      end
      if(flush) begin
        write_ptr <= 3'b000;
      end else begin
        if(ports_s_ports_fire) begin
          write_ptr <= (write_ptr + 3'b001);
        end
      end
      if(flush) begin
        fifo_cnt <= 3'b000;
      end else begin
        if(when_FIFO_l61) begin
          fifo_cnt <= (fifo_cnt + 3'b001);
        end else begin
          if(when_FIFO_l64) begin
            fifo_cnt <= (fifo_cnt - 3'b001);
          end
        end
      end
    end
  end

  always @(posedge io_axiClk) begin
    if(!flush) begin
      if(ports_s_ports_fire) begin
        if(_zz_1[0]) begin
          fifo_ram_0 <= ports_s_ports_payload;
        end
        if(_zz_1[1]) begin
          fifo_ram_1 <= ports_s_ports_payload;
        end
        if(_zz_1[2]) begin
          fifo_ram_2 <= ports_s_ports_payload;
        end
        if(_zz_1[3]) begin
          fifo_ram_3 <= ports_s_ports_payload;
        end
      end
    end
  end


endmodule

module StreamFifo (
  input               io_push_valid,
  output              io_push_ready,
  input               io_push_payload,
  output              io_pop_valid,
  input               io_pop_ready,
  output              io_pop_payload,
  input               io_flush,
  output     [1:0]    io_occupancy,
  output     [1:0]    io_availability,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  reg        [0:0]    _zz_logic_ram_port0;
  wire                _zz_logic_ram_port;
  wire                _zz_io_pop_payload;
  wire       [0:0]    _zz_logic_ram_port_1;
  wire       [0:0]    _zz_io_availability;
  reg                 _zz_1;
  reg                 logic_pushPtr_willIncrement;
  reg                 logic_pushPtr_willClear;
  reg        [0:0]    logic_pushPtr_valueNext;
  reg        [0:0]    logic_pushPtr_value;
  wire                logic_pushPtr_willOverflowIfInc;
  wire                logic_pushPtr_willOverflow;
  reg                 logic_popPtr_willIncrement;
  reg                 logic_popPtr_willClear;
  reg        [0:0]    logic_popPtr_valueNext;
  reg        [0:0]    logic_popPtr_value;
  wire                logic_popPtr_willOverflowIfInc;
  wire                logic_popPtr_willOverflow;
  wire                logic_ptrMatch;
  reg                 logic_risingOccupancy;
  wire                logic_pushing;
  wire                logic_popping;
  wire                logic_empty;
  wire                logic_full;
  reg                 _zz_io_pop_valid;
  wire                when_Stream_l1122;
  wire       [0:0]    logic_ptrDif;
  reg [0:0] logic_ram [0:1];

  assign _zz_io_availability = (logic_popPtr_value - logic_pushPtr_value);
  assign _zz_io_pop_payload = 1'b1;
  assign _zz_logic_ram_port_1 = io_push_payload;
  always @(posedge io_axiClk) begin
    if(_zz_io_pop_payload) begin
      _zz_logic_ram_port0 <= logic_ram[logic_popPtr_valueNext];
    end
  end

  always @(posedge io_axiClk) begin
    if(_zz_1) begin
      logic_ram[logic_pushPtr_value] <= _zz_logic_ram_port_1;
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_pushing) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willIncrement = 1'b0;
    if(logic_pushing) begin
      logic_pushPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_pushPtr_willClear = 1'b1;
    end
  end

  assign logic_pushPtr_willOverflowIfInc = (logic_pushPtr_value == 1'b1);
  assign logic_pushPtr_willOverflow = (logic_pushPtr_willOverflowIfInc && logic_pushPtr_willIncrement);
  always @(*) begin
    logic_pushPtr_valueNext = (logic_pushPtr_value + logic_pushPtr_willIncrement);
    if(logic_pushPtr_willClear) begin
      logic_pushPtr_valueNext = 1'b0;
    end
  end

  always @(*) begin
    logic_popPtr_willIncrement = 1'b0;
    if(logic_popping) begin
      logic_popPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_popPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_popPtr_willClear = 1'b1;
    end
  end

  assign logic_popPtr_willOverflowIfInc = (logic_popPtr_value == 1'b1);
  assign logic_popPtr_willOverflow = (logic_popPtr_willOverflowIfInc && logic_popPtr_willIncrement);
  always @(*) begin
    logic_popPtr_valueNext = (logic_popPtr_value + logic_popPtr_willIncrement);
    if(logic_popPtr_willClear) begin
      logic_popPtr_valueNext = 1'b0;
    end
  end

  assign logic_ptrMatch = (logic_pushPtr_value == logic_popPtr_value);
  assign logic_pushing = (io_push_valid && io_push_ready);
  assign logic_popping = (io_pop_valid && io_pop_ready);
  assign logic_empty = (logic_ptrMatch && (! logic_risingOccupancy));
  assign logic_full = (logic_ptrMatch && logic_risingOccupancy);
  assign io_push_ready = (! logic_full);
  assign io_pop_valid = ((! logic_empty) && (! (_zz_io_pop_valid && (! logic_full))));
  assign io_pop_payload = _zz_logic_ram_port0[0];
  assign when_Stream_l1122 = (logic_pushing != logic_popping);
  assign logic_ptrDif = (logic_pushPtr_value - logic_popPtr_value);
  assign io_occupancy = {(logic_risingOccupancy && logic_ptrMatch),logic_ptrDif};
  assign io_availability = {((! logic_risingOccupancy) && logic_ptrMatch),_zz_io_availability};
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      logic_pushPtr_value <= 1'b0;
      logic_popPtr_value <= 1'b0;
      logic_risingOccupancy <= 1'b0;
      _zz_io_pop_valid <= 1'b0;
    end else begin
      logic_pushPtr_value <= logic_pushPtr_valueNext;
      logic_popPtr_value <= logic_popPtr_valueNext;
      _zz_io_pop_valid <= (logic_popPtr_valueNext == logic_pushPtr_value);
      if(when_Stream_l1122) begin
        logic_risingOccupancy <= logic_pushing;
      end
      if(io_flush) begin
        logic_risingOccupancy <= 1'b0;
      end
    end
  end


endmodule

module StreamTransactionExtender (
  input      [6:0]    io_count,
  input               io_input_valid,
  output              io_input_ready,
  input      [63:0]   io_input_payload_data,
  input      [7:0]    io_input_payload_strb,
  input               io_input_payload_last,
  output              io_output_valid,
  input               io_output_ready,
  output     [63:0]   io_output_payload_data,
  output     [7:0]    io_output_payload_strb,
  output              io_output_payload_last,
  output              io_working,
  output              io_first,
  output              io_last,
  output              io_done,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  wire                counter_io_available;
  wire                counter_io_working;
  wire                counter_io_last;
  wire                counter_io_done;
  wire       [6:0]    counter_io_value;
  wire                io_input_fire;
  wire                io_output_fire;
  reg        [63:0]   payloadReg_data;
  reg        [7:0]    payloadReg_strb;
  reg                 payloadReg_last;
  wire       [63:0]   payload_data;
  wire       [7:0]    payload_strb;
  wire                payload_last;
  wire                io_input_fire_1;

  StreamTransactionCounter_6 counter (
    .io_ctrlFire        (io_input_fire        ), //i
    .io_targetFire      (io_output_fire       ), //i
    .io_available       (counter_io_available ), //o
    .io_count           (io_count[6:0]        ), //i
    .io_working         (counter_io_working   ), //o
    .io_last            (counter_io_last      ), //o
    .io_done            (counter_io_done      ), //o
    .io_value           (counter_io_value[6:0]), //o
    .io_axiClk          (io_axiClk            ), //i
    .resetCtrl_axiReset (resetCtrl_axiReset   )  //i
  );
  assign io_input_fire = (io_input_valid && io_input_ready);
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign payload_data = payloadReg_data;
  assign payload_strb = payloadReg_strb;
  assign payload_last = payloadReg_last;
  assign io_input_fire_1 = (io_input_valid && io_input_ready);
  assign io_output_payload_data = payload_data;
  assign io_output_payload_strb = payload_strb;
  assign io_output_payload_last = (counter_io_last && payload_last);
  assign io_output_valid = counter_io_working;
  assign io_input_ready = counter_io_available;
  assign io_last = counter_io_last;
  assign io_done = counter_io_done;
  assign io_first = ((counter_io_value == 7'h0) && counter_io_working);
  assign io_working = counter_io_working;
  always @(posedge io_axiClk) begin
    if(io_input_fire_1) begin
      payloadReg_data <= io_input_payload_data;
      payloadReg_strb <= io_input_payload_strb;
      payloadReg_last <= io_input_payload_last;
    end
  end


endmodule

//StreamTransactionCounter_1 replaced by StreamTransactionCounter

module StreamTransactionCounter (
  input               io_ctrlFire,
  input               io_targetFire,
  output              io_available,
  input      [7:0]    io_count,
  output              io_working,
  output              io_last,
  output              io_done,
  output     [7:0]    io_value,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  wire       [7:0]    _zz_counter_valueNext;
  wire       [0:0]    _zz_counter_valueNext_1;
  reg        [7:0]    expected;
  reg        [7:0]    countReg;
  reg                 counter_willIncrement;
  reg                 counter_willClear;
  reg        [7:0]    counter_valueNext;
  reg        [7:0]    counter_value;
  wire                counter_willOverflowIfInc;
  wire                counter_willOverflow;
  wire                lastOne;
  reg                 running;
  reg                 working;
  wire                done;
  wire                when_Stream_l1891;

  assign _zz_counter_valueNext_1 = counter_willIncrement;
  assign _zz_counter_valueNext = {7'd0, _zz_counter_valueNext_1};
  always @(*) begin
    expected = countReg;
    if(io_ctrlFire) begin
      expected = io_count;
    end
  end

  always @(*) begin
    counter_willIncrement = 1'b0;
    if(!done) begin
      if(when_Stream_l1891) begin
        counter_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    counter_willClear = 1'b0;
    if(done) begin
      counter_willClear = 1'b1;
    end
  end

  assign counter_willOverflowIfInc = (counter_value == 8'hff);
  assign counter_willOverflow = (counter_willOverflowIfInc && counter_willIncrement);
  always @(*) begin
    counter_valueNext = (counter_value + _zz_counter_valueNext);
    if(counter_willClear) begin
      counter_valueNext = 8'h0;
    end
  end

  assign lastOne = (expected <= counter_value);
  always @(*) begin
    working = running;
    if(io_ctrlFire) begin
      working = 1'b1;
    end
  end

  assign done = (lastOne && io_targetFire);
  assign when_Stream_l1891 = (io_targetFire && working);
  assign io_working = working;
  assign io_last = (lastOne && working);
  assign io_done = (done && working);
  assign io_value = counter_value;
  assign io_available = (! running);
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      counter_value <= 8'h0;
      running <= 1'b0;
    end else begin
      counter_value <= counter_valueNext;
      if(done) begin
        running <= 1'b0;
      end else begin
        running <= working;
      end
    end
  end

  always @(posedge io_axiClk) begin
    countReg <= expected;
  end


endmodule

//Axi4DownsizerSubTransactionGenerator replaced by Axi4DownsizerSubTransactionGenerator_1

module StreamTransactionExtender_2 (
  input      [6:0]    io_count,
  input               io_input_valid,
  output              io_input_ready,
  input      [6:0]    io_input_payload_ratio,
  input      [2:0]    io_input_payload_size,
  input      [7:0]    io_input_payload_len,
  input      [31:0]   io_input_payload_start,
  output              io_output_valid,
  input               io_output_ready,
  output     [6:0]    io_output_payload_ratio,
  output     [2:0]    io_output_payload_size,
  output     [7:0]    io_output_payload_len,
  output     [31:0]   io_output_payload_start,
  output              io_working,
  output              io_first,
  output              io_last,
  output              io_done,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  wire                counter_io_available;
  wire                counter_io_working;
  wire                counter_io_last;
  wire                counter_io_done;
  wire       [6:0]    counter_io_value;
  wire                io_input_fire;
  wire                io_output_fire;
  reg        [6:0]    payloadReg_ratio;
  reg        [2:0]    payloadReg_size;
  reg        [7:0]    payloadReg_len;
  reg        [31:0]   payloadReg_start;
  wire       [6:0]    payload_ratio;
  wire       [2:0]    payload_size;
  wire       [7:0]    payload_len;
  wire       [31:0]   payload_start;
  wire                io_input_fire_1;

  StreamTransactionCounter_6 counter (
    .io_ctrlFire        (io_input_fire        ), //i
    .io_targetFire      (io_output_fire       ), //i
    .io_available       (counter_io_available ), //o
    .io_count           (io_count[6:0]        ), //i
    .io_working         (counter_io_working   ), //o
    .io_last            (counter_io_last      ), //o
    .io_done            (counter_io_done      ), //o
    .io_value           (counter_io_value[6:0]), //o
    .io_axiClk          (io_axiClk            ), //i
    .resetCtrl_axiReset (resetCtrl_axiReset   )  //i
  );
  assign io_input_fire = (io_input_valid && io_input_ready);
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign payload_ratio = payloadReg_ratio;
  assign payload_size = payloadReg_size;
  assign payload_len = payloadReg_len;
  assign payload_start = payloadReg_start;
  assign io_input_fire_1 = (io_input_valid && io_input_ready);
  assign io_output_payload_ratio = payload_ratio;
  assign io_output_payload_size = payload_size;
  assign io_output_payload_len = payload_len;
  assign io_output_payload_start = payload_start;
  assign io_output_valid = counter_io_working;
  assign io_input_ready = counter_io_available;
  assign io_last = counter_io_last;
  assign io_done = counter_io_done;
  assign io_first = ((counter_io_value == 7'h0) && counter_io_working);
  assign io_working = counter_io_working;
  always @(posedge io_axiClk) begin
    if(io_input_fire_1) begin
      payloadReg_ratio <= io_input_payload_ratio;
      payloadReg_size <= io_input_payload_size;
      payloadReg_len <= io_input_payload_len;
      payloadReg_start <= io_input_payload_start;
    end
  end


endmodule

module StreamTransactionExtender_1 (
  input      [7:0]    io_count,
  input               io_input_valid,
  output              io_input_ready,
  input      [6:0]    io_input_payload_ratio,
  input      [2:0]    io_input_payload_size,
  input      [7:0]    io_input_payload_len,
  input      [31:0]   io_input_payload_start,
  output              io_output_valid,
  input               io_output_ready,
  output     [6:0]    io_output_payload_ratio,
  output     [2:0]    io_output_payload_size,
  output     [7:0]    io_output_payload_len,
  output     [31:0]   io_output_payload_start,
  output              io_working,
  output              io_first,
  output              io_last,
  output              io_done,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  wire                counter_io_available;
  wire                counter_io_working;
  wire                counter_io_last;
  wire                counter_io_done;
  wire       [7:0]    counter_io_value;
  wire                io_input_fire;
  wire                io_output_fire;
  reg        [6:0]    payloadReg_ratio;
  reg        [2:0]    payloadReg_size;
  reg        [7:0]    payloadReg_len;
  reg        [31:0]   payloadReg_start;
  wire       [6:0]    payload_ratio;
  wire       [2:0]    payload_size;
  wire       [7:0]    payload_len;
  wire       [31:0]   payload_start;
  wire                io_input_fire_1;

  StreamTransactionCounter_4 counter (
    .io_ctrlFire        (io_input_fire        ), //i
    .io_targetFire      (io_output_fire       ), //i
    .io_available       (counter_io_available ), //o
    .io_count           (io_count[7:0]        ), //i
    .io_working         (counter_io_working   ), //o
    .io_last            (counter_io_last      ), //o
    .io_done            (counter_io_done      ), //o
    .io_value           (counter_io_value[7:0]), //o
    .io_axiClk          (io_axiClk            ), //i
    .resetCtrl_axiReset (resetCtrl_axiReset   )  //i
  );
  assign io_input_fire = (io_input_valid && io_input_ready);
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign payload_ratio = payloadReg_ratio;
  assign payload_size = payloadReg_size;
  assign payload_len = payloadReg_len;
  assign payload_start = payloadReg_start;
  assign io_input_fire_1 = (io_input_valid && io_input_ready);
  assign io_output_payload_ratio = payload_ratio;
  assign io_output_payload_size = payload_size;
  assign io_output_payload_len = payload_len;
  assign io_output_payload_start = payload_start;
  assign io_output_valid = counter_io_working;
  assign io_input_ready = counter_io_available;
  assign io_last = counter_io_last;
  assign io_done = counter_io_done;
  assign io_first = ((counter_io_value == 8'h0) && counter_io_working);
  assign io_working = counter_io_working;
  always @(posedge io_axiClk) begin
    if(io_input_fire_1) begin
      payloadReg_ratio <= io_input_payload_ratio;
      payloadReg_size <= io_input_payload_size;
      payloadReg_len <= io_input_payload_len;
      payloadReg_start <= io_input_payload_start;
    end
  end


endmodule

module Axi4DownsizerSubTransactionGenerator_1 (
  input               io_input_valid,
  output              io_input_ready,
  input      [31:0]   io_input_payload_addr,
  input      [3:0]    io_input_payload_id,
  input      [3:0]    io_input_payload_region,
  input      [7:0]    io_input_payload_len,
  input      [2:0]    io_input_payload_size,
  input      [1:0]    io_input_payload_burst,
  input      [0:0]    io_input_payload_lock,
  input      [3:0]    io_input_payload_cache,
  input      [3:0]    io_input_payload_qos,
  input      [2:0]    io_input_payload_prot,
  output              io_output_valid,
  input               io_output_ready,
  output     [31:0]   io_output_payload_addr,
  output     [3:0]    io_output_payload_id,
  output     [3:0]    io_output_payload_region,
  output     [7:0]    io_output_payload_len,
  output     [2:0]    io_output_payload_size,
  output     [1:0]    io_output_payload_burst,
  output     [0:0]    io_output_payload_lock,
  output     [3:0]    io_output_payload_cache,
  output     [3:0]    io_output_payload_qos,
  output     [2:0]    io_output_payload_prot,
  output     [31:0]   io_start,
  output reg [6:0]    io_ratio,
  output reg [2:0]    io_size,
  output              io_working,
  output              io_last,
  output              io_done,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  wire                cmdExtender_io_input_ready;
  wire                cmdExtender_io_output_valid;
  wire       [31:0]   cmdExtender_io_output_payload_addr;
  wire       [3:0]    cmdExtender_io_output_payload_id;
  wire       [3:0]    cmdExtender_io_output_payload_region;
  wire       [7:0]    cmdExtender_io_output_payload_len;
  wire       [2:0]    cmdExtender_io_output_payload_size;
  wire       [1:0]    cmdExtender_io_output_payload_burst;
  wire       [0:0]    cmdExtender_io_output_payload_lock;
  wire       [3:0]    cmdExtender_io_output_payload_cache;
  wire       [3:0]    cmdExtender_io_output_payload_qos;
  wire       [2:0]    cmdExtender_io_output_payload_prot;
  wire                cmdExtender_io_working;
  wire                cmdExtender_io_first;
  wire                cmdExtender_io_last;
  wire                cmdExtender_io_done;
  wire       [31:0]   _zz_startAddress;
  wire       [6:0]    _zz_ratio;
  wire       [31:0]   _zz_address;
  wire       [15:0]   _zz_address_1;
  wire       [8:0]    _zz_address_2;
  wire       [8:0]    _zz_address_3;
  wire       [1:0]    _zz_address_4;
  reg        [31:0]   startAddress;
  wire       [2:0]    sizeDiff;
  reg        [2:0]    sizePerTrans;
  reg        [6:0]    ratio;
  wire                when_Axi4Downsizer_l45;
  wire                cmdStreamWithSize_valid;
  wire                cmdStreamWithSize_ready;
  wire       [31:0]   cmdStreamWithSize_payload_addr;
  wire       [3:0]    cmdStreamWithSize_payload_id;
  wire       [3:0]    cmdStreamWithSize_payload_region;
  wire       [7:0]    cmdStreamWithSize_payload_len;
  wire       [2:0]    cmdStreamWithSize_payload_size;
  wire       [1:0]    cmdStreamWithSize_payload_burst;
  wire       [0:0]    cmdStreamWithSize_payload_lock;
  wire       [3:0]    cmdStreamWithSize_payload_cache;
  wire       [3:0]    cmdStreamWithSize_payload_qos;
  wire       [2:0]    cmdStreamWithSize_payload_prot;
  wire                io_input_fire;
  reg        [2:0]    size;
  wire                cmdExtendedStream_valid;
  wire                cmdExtendedStream_ready;
  wire       [31:0]   cmdExtendedStream_payload_addr;
  wire       [3:0]    cmdExtendedStream_payload_id;
  wire       [3:0]    cmdExtendedStream_payload_region;
  wire       [7:0]    cmdExtendedStream_payload_len;
  wire       [2:0]    cmdExtendedStream_payload_size;
  wire       [1:0]    cmdExtendedStream_payload_burst;
  wire       [0:0]    cmdExtendedStream_payload_lock;
  wire       [3:0]    cmdExtendedStream_payload_cache;
  wire       [3:0]    cmdExtendedStream_payload_qos;
  wire       [2:0]    cmdExtendedStream_payload_prot;
  reg        [31:0]   address;
  wire                cmdStreamWithSize_fire;
  wire                cmdExtendedStream_fire;
  wire                cmdStream_valid;
  wire                cmdStream_ready;
  wire       [31:0]   cmdStream_payload_addr;
  wire       [3:0]    cmdStream_payload_id;
  wire       [3:0]    cmdStream_payload_region;
  wire       [7:0]    cmdStream_payload_len;
  wire       [2:0]    cmdStream_payload_size;
  wire       [1:0]    cmdStream_payload_burst;
  wire       [0:0]    cmdStream_payload_lock;
  wire       [3:0]    cmdStream_payload_cache;
  wire       [3:0]    cmdStream_payload_qos;
  wire       [2:0]    cmdStream_payload_prot;
  wire                io_input_fire_1;
  reg        [6:0]    dataRatio;
  wire                io_input_fire_2;

  assign _zz_startAddress = (io_input_payload_addr >>> io_input_payload_size);
  assign _zz_ratio = (7'h01 <<< sizeDiff);
  assign _zz_address_1 = ({7'd0,_zz_address_2} <<< size);
  assign _zz_address = {16'd0, _zz_address_1};
  assign _zz_address_2 = ({1'b0,cmdExtendedStream_payload_len} + _zz_address_3);
  assign _zz_address_4 = {1'b0,1'b1};
  assign _zz_address_3 = {7'd0, _zz_address_4};
  StreamTransactionExtender_4 cmdExtender (
    .io_count                 (ratio[6:0]                               ), //i
    .io_input_valid           (cmdStreamWithSize_valid                  ), //i
    .io_input_ready           (cmdExtender_io_input_ready               ), //o
    .io_input_payload_addr    (cmdStreamWithSize_payload_addr[31:0]     ), //i
    .io_input_payload_id      (cmdStreamWithSize_payload_id[3:0]        ), //i
    .io_input_payload_region  (cmdStreamWithSize_payload_region[3:0]    ), //i
    .io_input_payload_len     (cmdStreamWithSize_payload_len[7:0]       ), //i
    .io_input_payload_size    (cmdStreamWithSize_payload_size[2:0]      ), //i
    .io_input_payload_burst   (cmdStreamWithSize_payload_burst[1:0]     ), //i
    .io_input_payload_lock    (cmdStreamWithSize_payload_lock           ), //i
    .io_input_payload_cache   (cmdStreamWithSize_payload_cache[3:0]     ), //i
    .io_input_payload_qos     (cmdStreamWithSize_payload_qos[3:0]       ), //i
    .io_input_payload_prot    (cmdStreamWithSize_payload_prot[2:0]      ), //i
    .io_output_valid          (cmdExtender_io_output_valid              ), //o
    .io_output_ready          (cmdExtendedStream_ready                  ), //i
    .io_output_payload_addr   (cmdExtender_io_output_payload_addr[31:0] ), //o
    .io_output_payload_id     (cmdExtender_io_output_payload_id[3:0]    ), //o
    .io_output_payload_region (cmdExtender_io_output_payload_region[3:0]), //o
    .io_output_payload_len    (cmdExtender_io_output_payload_len[7:0]   ), //o
    .io_output_payload_size   (cmdExtender_io_output_payload_size[2:0]  ), //o
    .io_output_payload_burst  (cmdExtender_io_output_payload_burst[1:0] ), //o
    .io_output_payload_lock   (cmdExtender_io_output_payload_lock       ), //o
    .io_output_payload_cache  (cmdExtender_io_output_payload_cache[3:0] ), //o
    .io_output_payload_qos    (cmdExtender_io_output_payload_qos[3:0]   ), //o
    .io_output_payload_prot   (cmdExtender_io_output_payload_prot[2:0]  ), //o
    .io_working               (cmdExtender_io_working                   ), //o
    .io_first                 (cmdExtender_io_first                     ), //o
    .io_last                  (cmdExtender_io_last                      ), //o
    .io_done                  (cmdExtender_io_done                      ), //o
    .io_axiClk                (io_axiClk                                ), //i
    .resetCtrl_axiReset       (resetCtrl_axiReset                       )  //i
  );
  assign sizeDiff = (io_input_payload_size - 3'b010);
  assign when_Axi4Downsizer_l45 = (3'b010 < io_input_payload_size);
  always @(*) begin
    if(when_Axi4Downsizer_l45) begin
      startAddress = (_zz_startAddress <<< io_input_payload_size);
    end else begin
      startAddress = io_input_payload_addr;
    end
  end

  always @(*) begin
    if(when_Axi4Downsizer_l45) begin
      ratio = (_zz_ratio - 7'h01);
    end else begin
      ratio = 7'h0;
    end
  end

  always @(*) begin
    if(when_Axi4Downsizer_l45) begin
      sizePerTrans = 3'b010;
    end else begin
      sizePerTrans = io_input_payload_size;
    end
  end

  assign cmdStreamWithSize_valid = io_input_valid;
  assign io_input_ready = cmdStreamWithSize_ready;
  assign cmdStreamWithSize_payload_addr = startAddress;
  assign cmdStreamWithSize_payload_size = sizePerTrans;
  assign cmdStreamWithSize_payload_id = io_input_payload_id;
  assign cmdStreamWithSize_payload_region = io_input_payload_region;
  assign cmdStreamWithSize_payload_len = io_input_payload_len;
  assign cmdStreamWithSize_payload_burst = io_input_payload_burst;
  assign cmdStreamWithSize_payload_lock = io_input_payload_lock;
  assign cmdStreamWithSize_payload_cache = io_input_payload_cache;
  assign cmdStreamWithSize_payload_qos = io_input_payload_qos;
  assign cmdStreamWithSize_payload_prot = io_input_payload_prot;
  assign io_input_fire = (io_input_valid && io_input_ready);
  assign cmdStreamWithSize_ready = cmdExtender_io_input_ready;
  assign cmdExtendedStream_valid = cmdExtender_io_output_valid;
  assign cmdExtendedStream_payload_addr = cmdExtender_io_output_payload_addr;
  assign cmdExtendedStream_payload_id = cmdExtender_io_output_payload_id;
  assign cmdExtendedStream_payload_region = cmdExtender_io_output_payload_region;
  assign cmdExtendedStream_payload_len = cmdExtender_io_output_payload_len;
  assign cmdExtendedStream_payload_size = cmdExtender_io_output_payload_size;
  assign cmdExtendedStream_payload_burst = cmdExtender_io_output_payload_burst;
  assign cmdExtendedStream_payload_lock = cmdExtender_io_output_payload_lock;
  assign cmdExtendedStream_payload_cache = cmdExtender_io_output_payload_cache;
  assign cmdExtendedStream_payload_qos = cmdExtender_io_output_payload_qos;
  assign cmdExtendedStream_payload_prot = cmdExtender_io_output_payload_prot;
  assign cmdStreamWithSize_fire = (cmdStreamWithSize_valid && cmdStreamWithSize_ready);
  assign cmdExtendedStream_fire = (cmdExtendedStream_valid && cmdExtendedStream_ready);
  assign cmdStream_valid = cmdExtendedStream_valid;
  assign cmdExtendedStream_ready = cmdStream_ready;
  assign cmdStream_payload_addr = address;
  assign cmdStream_payload_id = cmdExtendedStream_payload_id;
  assign cmdStream_payload_region = cmdExtendedStream_payload_region;
  assign cmdStream_payload_len = cmdExtendedStream_payload_len;
  assign cmdStream_payload_size = cmdExtendedStream_payload_size;
  assign cmdStream_payload_burst = cmdExtendedStream_payload_burst;
  assign cmdStream_payload_lock = cmdExtendedStream_payload_lock;
  assign cmdStream_payload_cache = cmdExtendedStream_payload_cache;
  assign cmdStream_payload_qos = cmdExtendedStream_payload_qos;
  assign cmdStream_payload_prot = cmdExtendedStream_payload_prot;
  assign io_input_fire_1 = (io_input_valid && io_input_ready);
  assign io_input_fire_2 = (io_input_valid && io_input_ready);
  always @(*) begin
    if(io_input_fire_2) begin
      io_ratio = ratio;
    end else begin
      io_ratio = dataRatio;
    end
  end

  always @(*) begin
    if(io_input_fire_2) begin
      io_size = sizePerTrans;
    end else begin
      io_size = size;
    end
  end

  assign io_working = cmdExtender_io_working;
  assign io_last = cmdExtender_io_last;
  assign io_done = cmdExtender_io_done;
  assign io_start = startAddress;
  assign io_output_valid = cmdStream_valid;
  assign cmdStream_ready = io_output_ready;
  assign io_output_payload_addr = cmdStream_payload_addr;
  assign io_output_payload_id = cmdStream_payload_id;
  assign io_output_payload_region = cmdStream_payload_region;
  assign io_output_payload_len = cmdStream_payload_len;
  assign io_output_payload_size = cmdStream_payload_size;
  assign io_output_payload_burst = cmdStream_payload_burst;
  assign io_output_payload_lock = cmdStream_payload_lock;
  assign io_output_payload_cache = cmdStream_payload_cache;
  assign io_output_payload_qos = cmdStream_payload_qos;
  assign io_output_payload_prot = cmdStream_payload_prot;
  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      size <= 3'b010;
      address <= 32'h0;
      dataRatio <= 7'h0;
    end else begin
      if(io_input_fire) begin
        size <= sizePerTrans;
      end
      if(cmdStreamWithSize_fire) begin
        address <= cmdStreamWithSize_payload_addr;
      end else begin
        if(cmdExtendedStream_fire) begin
          address <= (address + _zz_address);
        end
      end
      if(io_input_fire_1) begin
        dataRatio <= ratio;
      end
    end
  end


endmodule

//StreamTransactionCounter_2 replaced by StreamTransactionCounter_6

//StreamTransactionExtender_3 replaced by StreamTransactionExtender_4

//StreamTransactionCounter_3 replaced by StreamTransactionCounter_6

module StreamTransactionCounter_4 (
  input               io_ctrlFire,
  input               io_targetFire,
  output              io_available,
  input      [7:0]    io_count,
  output              io_working,
  output              io_last,
  output              io_done,
  output     [7:0]    io_value,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  wire       [7:0]    _zz_counter_valueNext;
  wire       [0:0]    _zz_counter_valueNext_1;
  reg        [7:0]    countReg;
  reg                 counter_willIncrement;
  reg                 counter_willClear;
  reg        [7:0]    counter_valueNext;
  reg        [7:0]    counter_value;
  wire                counter_willOverflowIfInc;
  wire                counter_willOverflow;
  wire       [7:0]    expected;
  wire                lastOne;
  reg                 running;
  wire                working;
  wire                done;
  wire                when_Stream_l1891;

  assign _zz_counter_valueNext_1 = counter_willIncrement;
  assign _zz_counter_valueNext = {7'd0, _zz_counter_valueNext_1};
  always @(*) begin
    counter_willIncrement = 1'b0;
    if(!done) begin
      if(when_Stream_l1891) begin
        counter_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    counter_willClear = 1'b0;
    if(done) begin
      counter_willClear = 1'b1;
    end
  end

  assign counter_willOverflowIfInc = (counter_value == 8'hff);
  assign counter_willOverflow = (counter_willOverflowIfInc && counter_willIncrement);
  always @(*) begin
    counter_valueNext = (counter_value + _zz_counter_valueNext);
    if(counter_willClear) begin
      counter_valueNext = 8'h0;
    end
  end

  assign expected = countReg;
  assign lastOne = (expected <= counter_value);
  assign working = running;
  assign done = (lastOne && io_targetFire);
  assign when_Stream_l1891 = (io_targetFire && working);
  assign io_working = working;
  assign io_last = (lastOne && working);
  assign io_done = (done && working);
  assign io_value = counter_value;
  assign io_available = ((! working) || io_done);
  always @(posedge io_axiClk) begin
    if(io_ctrlFire) begin
      countReg <= io_count;
    end
  end

  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      counter_value <= 8'h0;
      running <= 1'b0;
    end else begin
      counter_value <= counter_valueNext;
      if(io_ctrlFire) begin
        running <= 1'b1;
      end else begin
        if(done) begin
          running <= 1'b0;
        end
      end
    end
  end


endmodule

module StreamTransactionExtender_4 (
  input      [6:0]    io_count,
  input               io_input_valid,
  output              io_input_ready,
  input      [31:0]   io_input_payload_addr,
  input      [3:0]    io_input_payload_id,
  input      [3:0]    io_input_payload_region,
  input      [7:0]    io_input_payload_len,
  input      [2:0]    io_input_payload_size,
  input      [1:0]    io_input_payload_burst,
  input      [0:0]    io_input_payload_lock,
  input      [3:0]    io_input_payload_cache,
  input      [3:0]    io_input_payload_qos,
  input      [2:0]    io_input_payload_prot,
  output              io_output_valid,
  input               io_output_ready,
  output     [31:0]   io_output_payload_addr,
  output     [3:0]    io_output_payload_id,
  output     [3:0]    io_output_payload_region,
  output     [7:0]    io_output_payload_len,
  output     [2:0]    io_output_payload_size,
  output     [1:0]    io_output_payload_burst,
  output     [0:0]    io_output_payload_lock,
  output     [3:0]    io_output_payload_cache,
  output     [3:0]    io_output_payload_qos,
  output     [2:0]    io_output_payload_prot,
  output              io_working,
  output              io_first,
  output              io_last,
  output              io_done,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  wire                counter_io_available;
  wire                counter_io_working;
  wire                counter_io_last;
  wire                counter_io_done;
  wire       [6:0]    counter_io_value;
  wire                io_input_fire;
  wire                io_output_fire;
  reg        [31:0]   payloadReg_addr;
  reg        [3:0]    payloadReg_id;
  reg        [3:0]    payloadReg_region;
  reg        [7:0]    payloadReg_len;
  reg        [2:0]    payloadReg_size;
  reg        [1:0]    payloadReg_burst;
  reg        [0:0]    payloadReg_lock;
  reg        [3:0]    payloadReg_cache;
  reg        [3:0]    payloadReg_qos;
  reg        [2:0]    payloadReg_prot;
  wire       [31:0]   payload_addr;
  wire       [3:0]    payload_id;
  wire       [3:0]    payload_region;
  wire       [7:0]    payload_len;
  wire       [2:0]    payload_size;
  wire       [1:0]    payload_burst;
  wire       [0:0]    payload_lock;
  wire       [3:0]    payload_cache;
  wire       [3:0]    payload_qos;
  wire       [2:0]    payload_prot;
  wire                io_input_fire_1;

  StreamTransactionCounter_6 counter (
    .io_ctrlFire        (io_input_fire        ), //i
    .io_targetFire      (io_output_fire       ), //i
    .io_available       (counter_io_available ), //o
    .io_count           (io_count[6:0]        ), //i
    .io_working         (counter_io_working   ), //o
    .io_last            (counter_io_last      ), //o
    .io_done            (counter_io_done      ), //o
    .io_value           (counter_io_value[6:0]), //o
    .io_axiClk          (io_axiClk            ), //i
    .resetCtrl_axiReset (resetCtrl_axiReset   )  //i
  );
  assign io_input_fire = (io_input_valid && io_input_ready);
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign payload_addr = payloadReg_addr;
  assign payload_id = payloadReg_id;
  assign payload_region = payloadReg_region;
  assign payload_len = payloadReg_len;
  assign payload_size = payloadReg_size;
  assign payload_burst = payloadReg_burst;
  assign payload_lock = payloadReg_lock;
  assign payload_cache = payloadReg_cache;
  assign payload_qos = payloadReg_qos;
  assign payload_prot = payloadReg_prot;
  assign io_input_fire_1 = (io_input_valid && io_input_ready);
  assign io_output_payload_addr = payload_addr;
  assign io_output_payload_id = payload_id;
  assign io_output_payload_region = payload_region;
  assign io_output_payload_len = payload_len;
  assign io_output_payload_size = payload_size;
  assign io_output_payload_burst = payload_burst;
  assign io_output_payload_lock = payload_lock;
  assign io_output_payload_cache = payload_cache;
  assign io_output_payload_qos = payload_qos;
  assign io_output_payload_prot = payload_prot;
  assign io_output_valid = counter_io_working;
  assign io_input_ready = counter_io_available;
  assign io_last = counter_io_last;
  assign io_done = counter_io_done;
  assign io_first = ((counter_io_value == 7'h0) && counter_io_working);
  assign io_working = counter_io_working;
  always @(posedge io_axiClk) begin
    if(io_input_fire_1) begin
      payloadReg_addr <= io_input_payload_addr;
      payloadReg_id <= io_input_payload_id;
      payloadReg_region <= io_input_payload_region;
      payloadReg_len <= io_input_payload_len;
      payloadReg_size <= io_input_payload_size;
      payloadReg_burst <= io_input_payload_burst;
      payloadReg_lock <= io_input_payload_lock;
      payloadReg_cache <= io_input_payload_cache;
      payloadReg_qos <= io_input_payload_qos;
      payloadReg_prot <= io_input_payload_prot;
    end
  end


endmodule

//StreamTransactionCounter_5 replaced by StreamTransactionCounter_6

module StreamTransactionCounter_6 (
  input               io_ctrlFire,
  input               io_targetFire,
  output              io_available,
  input      [6:0]    io_count,
  output              io_working,
  output              io_last,
  output              io_done,
  output     [6:0]    io_value,
  input               io_axiClk,
  input               resetCtrl_axiReset
);

  wire       [6:0]    _zz_counter_valueNext;
  wire       [0:0]    _zz_counter_valueNext_1;
  reg        [6:0]    countReg;
  reg                 counter_willIncrement;
  reg                 counter_willClear;
  reg        [6:0]    counter_valueNext;
  reg        [6:0]    counter_value;
  wire                counter_willOverflowIfInc;
  wire                counter_willOverflow;
  wire       [6:0]    expected;
  wire                lastOne;
  reg                 running;
  wire                working;
  wire                done;
  wire                when_Stream_l1891;

  assign _zz_counter_valueNext_1 = counter_willIncrement;
  assign _zz_counter_valueNext = {6'd0, _zz_counter_valueNext_1};
  always @(*) begin
    counter_willIncrement = 1'b0;
    if(!done) begin
      if(when_Stream_l1891) begin
        counter_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    counter_willClear = 1'b0;
    if(done) begin
      counter_willClear = 1'b1;
    end
  end

  assign counter_willOverflowIfInc = (counter_value == 7'h7f);
  assign counter_willOverflow = (counter_willOverflowIfInc && counter_willIncrement);
  always @(*) begin
    counter_valueNext = (counter_value + _zz_counter_valueNext);
    if(counter_willClear) begin
      counter_valueNext = 7'h0;
    end
  end

  assign expected = countReg;
  assign lastOne = (expected <= counter_value);
  assign working = running;
  assign done = (lastOne && io_targetFire);
  assign when_Stream_l1891 = (io_targetFire && working);
  assign io_working = working;
  assign io_last = (lastOne && working);
  assign io_done = (done && working);
  assign io_value = counter_value;
  assign io_available = ((! working) || io_done);
  always @(posedge io_axiClk) begin
    if(io_ctrlFire) begin
      countReg <= io_count;
    end
  end

  always @(posedge io_axiClk or posedge resetCtrl_axiReset) begin
    if(resetCtrl_axiReset) begin
      counter_value <= 7'h0;
      running <= 1'b0;
    end else begin
      counter_value <= counter_valueNext;
      if(io_ctrlFire) begin
        running <= 1'b1;
      end else begin
        if(done) begin
          running <= 1'b0;
        end
      end
    end
  end


endmodule
