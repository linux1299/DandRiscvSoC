// Generator : SpinalHDL v1.8.1    git head : 2a7592004363e5b40ec43e1f122ed8641cd8965b
// Component : DandRiscvSimple
// Git hash  : 2642408e20774ae356a7923571e5e25dc672b2ab

`timescale 1ns/1ps

module DandRiscvSimple (
  output              icache_ar_valid,
  input               icache_ar_ready,
  output     [63:0]   icache_ar_payload_addr,
  output     [3:0]    icache_ar_payload_id,
  output     [7:0]    icache_ar_payload_len,
  output     [2:0]    icache_ar_payload_size,
  output     [1:0]    icache_ar_payload_burst,
  input               icache_r_valid,
  output              icache_r_ready,
  input      [63:0]   icache_r_payload_data,
  input      [3:0]    icache_r_payload_id,
  input      [1:0]    icache_r_payload_resp,
  input               icache_r_payload_last,
  output reg          dcache_ar_valid,
  input               dcache_ar_ready,
  output reg [63:0]   dcache_ar_payload_addr,
  output reg [3:0]    dcache_ar_payload_id,
  output reg [7:0]    dcache_ar_payload_len,
  output reg [2:0]    dcache_ar_payload_size,
  output reg [1:0]    dcache_ar_payload_burst,
  input               dcache_r_valid,
  output              dcache_r_ready,
  input      [63:0]   dcache_r_payload_data,
  input      [3:0]    dcache_r_payload_id,
  input      [1:0]    dcache_r_payload_resp,
  input               dcache_r_payload_last,
  output reg          dcache_aw_valid,
  input               dcache_aw_ready,
  output reg [63:0]   dcache_aw_payload_addr,
  output reg [3:0]    dcache_aw_payload_id,
  output reg [7:0]    dcache_aw_payload_len,
  output reg [2:0]    dcache_aw_payload_size,
  output reg [1:0]    dcache_aw_payload_burst,
  output reg          dcache_w_valid,
  input               dcache_w_ready,
  output reg [63:0]   dcache_w_payload_data,
  output reg [7:0]    dcache_w_payload_strb,
  output reg          dcache_w_payload_last,
  input               dcache_b_valid,
  output              dcache_b_ready,
  input      [3:0]    dcache_b_payload_id,
  input      [1:0]    dcache_b_payload_resp,
  input               clk,
  input               reset
);
  localparam CsrCtrlEnum_IDLE = 4'd0;
  localparam CsrCtrlEnum_ECALL = 4'd1;
  localparam CsrCtrlEnum_EBREAK = 4'd2;
  localparam CsrCtrlEnum_MRET = 4'd3;
  localparam CsrCtrlEnum_CSRRW = 4'd4;
  localparam CsrCtrlEnum_CSRRS = 4'd5;
  localparam CsrCtrlEnum_CSRRC = 4'd6;
  localparam CsrCtrlEnum_CSRRWI = 4'd7;
  localparam CsrCtrlEnum_CSRRSI = 4'd8;
  localparam CsrCtrlEnum_CSRRCI = 4'd9;
  localparam AluCtrlEnum_IDLE = 5'd0;
  localparam AluCtrlEnum_ADD = 5'd1;
  localparam AluCtrlEnum_SUB = 5'd2;
  localparam AluCtrlEnum_SLT = 5'd3;
  localparam AluCtrlEnum_SLTU = 5'd4;
  localparam AluCtrlEnum_XOR_1 = 5'd5;
  localparam AluCtrlEnum_SLL_1 = 5'd6;
  localparam AluCtrlEnum_SRL_1 = 5'd7;
  localparam AluCtrlEnum_SRA_1 = 5'd8;
  localparam AluCtrlEnum_AND_1 = 5'd9;
  localparam AluCtrlEnum_OR_1 = 5'd10;
  localparam AluCtrlEnum_LUI = 5'd11;
  localparam AluCtrlEnum_AUIPC = 5'd12;
  localparam AluCtrlEnum_JAL = 5'd13;
  localparam AluCtrlEnum_JALR = 5'd14;
  localparam AluCtrlEnum_BEQ = 5'd15;
  localparam AluCtrlEnum_BNE = 5'd16;
  localparam AluCtrlEnum_BLT = 5'd17;
  localparam AluCtrlEnum_BGE = 5'd18;
  localparam AluCtrlEnum_BLTU = 5'd19;
  localparam AluCtrlEnum_BGEU = 5'd20;
  localparam AluCtrlEnum_CSR = 5'd21;
  localparam MemCtrlEnum_IDLE = 4'd0;
  localparam MemCtrlEnum_LB = 4'd1;
  localparam MemCtrlEnum_LBU = 4'd2;
  localparam MemCtrlEnum_LH = 4'd3;
  localparam MemCtrlEnum_LHU = 4'd4;
  localparam MemCtrlEnum_LW = 4'd5;
  localparam MemCtrlEnum_LWU = 4'd6;
  localparam MemCtrlEnum_LD = 4'd7;
  localparam MemCtrlEnum_SB = 4'd8;
  localparam MemCtrlEnum_SH = 4'd9;
  localparam MemCtrlEnum_SW = 4'd10;
  localparam MemCtrlEnum_SD = 4'd11;

  wire                regFileModule_1_write_ports_rd_wen;
  wire                clint_1_ecall;
  wire                clint_1_ebreak;
  wire                clint_1_mret;
  wire       [63:0]   timer_1_addr;
  wire                iCache_1_sram_4_ports_rsp_valid;
  wire       [511:0]  iCache_1_sram_4_ports_rsp_payload_data;
  wire                iCache_1_sram_5_ports_rsp_valid;
  wire       [511:0]  iCache_1_sram_5_ports_rsp_payload_data;
  wire                iCache_1_sram_6_ports_rsp_valid;
  wire       [511:0]  iCache_1_sram_6_ports_rsp_payload_data;
  wire                iCache_1_sram_7_ports_rsp_valid;
  wire       [511:0]  iCache_1_sram_7_ports_rsp_payload_data;
  wire                iCache_1_sram_8_ports_rsp_valid;
  wire       [511:0]  iCache_1_sram_8_ports_rsp_payload_data;
  wire                iCache_1_sram_9_ports_rsp_valid;
  wire       [511:0]  iCache_1_sram_9_ports_rsp_payload_data;
  wire                iCache_1_sram_10_ports_rsp_valid;
  wire       [511:0]  iCache_1_sram_10_ports_rsp_payload_data;
  wire                iCache_1_sram_11_ports_rsp_valid;
  wire       [511:0]  iCache_1_sram_11_ports_rsp_payload_data;
  wire                iCache_1_sram_12_ports_rsp_valid;
  wire       [511:0]  iCache_1_sram_12_ports_rsp_payload_data;
  wire                iCache_1_sram_13_ports_rsp_valid;
  wire       [511:0]  iCache_1_sram_13_ports_rsp_payload_data;
  wire                iCache_1_sram_14_ports_rsp_valid;
  wire       [511:0]  iCache_1_sram_14_ports_rsp_payload_data;
  wire                iCache_1_sram_15_ports_rsp_valid;
  wire       [511:0]  iCache_1_sram_15_ports_rsp_payload_data;
  wire                dCache_1_next_level_cmd_ready;
  wire                dCache_1_next_level_rsp_valid;
  wire                fetch_FetchPlugin_pc_stream_fifo_ports_m_ports_valid;
  wire       [63:0]   fetch_FetchPlugin_pc_stream_fifo_ports_m_ports_payload;
  wire                fetch_FetchPlugin_pc_stream_fifo_ports_s_ports_ready;
  wire       [63:0]   fetch_FetchPlugin_pc_stream_fifo_next_payload;
  wire                fetch_FetchPlugin_pc_stream_fifo_next_valid;
  wire                fetch_FetchPlugin_predict_taken_fifo_ports_m_ports_valid;
  wire                fetch_FetchPlugin_predict_taken_fifo_ports_m_ports_payload;
  wire                fetch_FetchPlugin_predict_taken_fifo_ports_s_ports_ready;
  wire                fetch_FetchPlugin_instruction_stream_fifo_ports_m_ports_valid;
  wire       [31:0]   fetch_FetchPlugin_instruction_stream_fifo_ports_m_ports_payload;
  wire                fetch_FetchPlugin_instruction_stream_fifo_ports_s_ports_ready;
  wire                gshare_predictor_1_predict_taken;
  wire       [6:0]    gshare_predictor_1_predict_history;
  wire       [63:0]   gshare_predictor_1_predict_pc_next;
  wire       [63:0]   regFileModule_1_read_ports_rs1_value;
  wire       [63:0]   regFileModule_1_read_ports_rs2_value;
  wire       [63:0]   csrRegfile_1_cpu_ports_rdata;
  wire       [63:0]   csrRegfile_1_clint_ports_mtvec;
  wire       [63:0]   csrRegfile_1_clint_ports_mepc;
  wire       [63:0]   csrRegfile_1_clint_ports_mstatus;
  wire                csrRegfile_1_clint_ports_global_int_en;
  wire                csrRegfile_1_clint_ports_mtime_int_en;
  wire                csrRegfile_1_clint_ports_mtime_int_pend;
  wire                clint_1_csr_ports_mepc_wen;
  wire       [63:0]   clint_1_csr_ports_mepc_wdata;
  wire                clint_1_csr_ports_mcause_wen;
  wire       [63:0]   clint_1_csr_ports_mcause_wdata;
  wire                clint_1_csr_ports_mstatus_wen;
  wire       [63:0]   clint_1_csr_ports_mstatus_wdata;
  wire                clint_1_int_en;
  wire       [63:0]   clint_1_int_pc;
  wire                clint_1_int_hold;
  wire       [63:0]   timer_1_rdata;
  wire                timer_1_timer_int;
  wire                iCache_1_cpu_cmd_ready;
  wire                iCache_1_cpu_rsp_valid;
  wire       [31:0]   iCache_1_cpu_rsp_payload_data;
  wire                iCache_1_sram_0_ports_cmd_valid;
  wire       [6:0]    iCache_1_sram_0_ports_cmd_payload_addr;
  wire       [15:0]   iCache_1_sram_0_ports_cmd_payload_wen;
  wire       [511:0]  iCache_1_sram_0_ports_cmd_payload_wdata;
  wire       [63:0]   iCache_1_sram_0_ports_cmd_payload_wstrb;
  wire                iCache_1_sram_1_ports_cmd_valid;
  wire       [6:0]    iCache_1_sram_1_ports_cmd_payload_addr;
  wire       [15:0]   iCache_1_sram_1_ports_cmd_payload_wen;
  wire       [511:0]  iCache_1_sram_1_ports_cmd_payload_wdata;
  wire       [63:0]   iCache_1_sram_1_ports_cmd_payload_wstrb;
  wire                iCache_1_sram_2_ports_cmd_valid;
  wire       [6:0]    iCache_1_sram_2_ports_cmd_payload_addr;
  wire       [15:0]   iCache_1_sram_2_ports_cmd_payload_wen;
  wire       [511:0]  iCache_1_sram_2_ports_cmd_payload_wdata;
  wire       [63:0]   iCache_1_sram_2_ports_cmd_payload_wstrb;
  wire                iCache_1_sram_3_ports_cmd_valid;
  wire       [6:0]    iCache_1_sram_3_ports_cmd_payload_addr;
  wire       [15:0]   iCache_1_sram_3_ports_cmd_payload_wen;
  wire       [511:0]  iCache_1_sram_3_ports_cmd_payload_wdata;
  wire       [63:0]   iCache_1_sram_3_ports_cmd_payload_wstrb;
  wire                iCache_1_sram_4_ports_cmd_valid;
  wire       [6:0]    iCache_1_sram_4_ports_cmd_payload_addr;
  wire       [15:0]   iCache_1_sram_4_ports_cmd_payload_wen;
  wire       [511:0]  iCache_1_sram_4_ports_cmd_payload_wdata;
  wire       [63:0]   iCache_1_sram_4_ports_cmd_payload_wstrb;
  wire                iCache_1_sram_5_ports_cmd_valid;
  wire       [6:0]    iCache_1_sram_5_ports_cmd_payload_addr;
  wire       [15:0]   iCache_1_sram_5_ports_cmd_payload_wen;
  wire       [511:0]  iCache_1_sram_5_ports_cmd_payload_wdata;
  wire       [63:0]   iCache_1_sram_5_ports_cmd_payload_wstrb;
  wire                iCache_1_sram_6_ports_cmd_valid;
  wire       [6:0]    iCache_1_sram_6_ports_cmd_payload_addr;
  wire       [15:0]   iCache_1_sram_6_ports_cmd_payload_wen;
  wire       [511:0]  iCache_1_sram_6_ports_cmd_payload_wdata;
  wire       [63:0]   iCache_1_sram_6_ports_cmd_payload_wstrb;
  wire                iCache_1_sram_7_ports_cmd_valid;
  wire       [6:0]    iCache_1_sram_7_ports_cmd_payload_addr;
  wire       [15:0]   iCache_1_sram_7_ports_cmd_payload_wen;
  wire       [511:0]  iCache_1_sram_7_ports_cmd_payload_wdata;
  wire       [63:0]   iCache_1_sram_7_ports_cmd_payload_wstrb;
  wire                iCache_1_sram_8_ports_cmd_valid;
  wire       [6:0]    iCache_1_sram_8_ports_cmd_payload_addr;
  wire       [15:0]   iCache_1_sram_8_ports_cmd_payload_wen;
  wire       [511:0]  iCache_1_sram_8_ports_cmd_payload_wdata;
  wire       [63:0]   iCache_1_sram_8_ports_cmd_payload_wstrb;
  wire                iCache_1_sram_9_ports_cmd_valid;
  wire       [6:0]    iCache_1_sram_9_ports_cmd_payload_addr;
  wire       [15:0]   iCache_1_sram_9_ports_cmd_payload_wen;
  wire       [511:0]  iCache_1_sram_9_ports_cmd_payload_wdata;
  wire       [63:0]   iCache_1_sram_9_ports_cmd_payload_wstrb;
  wire                iCache_1_sram_10_ports_cmd_valid;
  wire       [6:0]    iCache_1_sram_10_ports_cmd_payload_addr;
  wire       [15:0]   iCache_1_sram_10_ports_cmd_payload_wen;
  wire       [511:0]  iCache_1_sram_10_ports_cmd_payload_wdata;
  wire       [63:0]   iCache_1_sram_10_ports_cmd_payload_wstrb;
  wire                iCache_1_sram_11_ports_cmd_valid;
  wire       [6:0]    iCache_1_sram_11_ports_cmd_payload_addr;
  wire       [15:0]   iCache_1_sram_11_ports_cmd_payload_wen;
  wire       [511:0]  iCache_1_sram_11_ports_cmd_payload_wdata;
  wire       [63:0]   iCache_1_sram_11_ports_cmd_payload_wstrb;
  wire                iCache_1_sram_12_ports_cmd_valid;
  wire       [6:0]    iCache_1_sram_12_ports_cmd_payload_addr;
  wire       [15:0]   iCache_1_sram_12_ports_cmd_payload_wen;
  wire       [511:0]  iCache_1_sram_12_ports_cmd_payload_wdata;
  wire       [63:0]   iCache_1_sram_12_ports_cmd_payload_wstrb;
  wire                iCache_1_sram_13_ports_cmd_valid;
  wire       [6:0]    iCache_1_sram_13_ports_cmd_payload_addr;
  wire       [15:0]   iCache_1_sram_13_ports_cmd_payload_wen;
  wire       [511:0]  iCache_1_sram_13_ports_cmd_payload_wdata;
  wire       [63:0]   iCache_1_sram_13_ports_cmd_payload_wstrb;
  wire                iCache_1_sram_14_ports_cmd_valid;
  wire       [6:0]    iCache_1_sram_14_ports_cmd_payload_addr;
  wire       [15:0]   iCache_1_sram_14_ports_cmd_payload_wen;
  wire       [511:0]  iCache_1_sram_14_ports_cmd_payload_wdata;
  wire       [63:0]   iCache_1_sram_14_ports_cmd_payload_wstrb;
  wire                iCache_1_sram_15_ports_cmd_valid;
  wire       [6:0]    iCache_1_sram_15_ports_cmd_payload_addr;
  wire       [15:0]   iCache_1_sram_15_ports_cmd_payload_wen;
  wire       [511:0]  iCache_1_sram_15_ports_cmd_payload_wdata;
  wire       [63:0]   iCache_1_sram_15_ports_cmd_payload_wstrb;
  wire                iCache_1_next_level_cmd_valid;
  wire       [63:0]   iCache_1_next_level_cmd_payload_addr;
  wire       [3:0]    iCache_1_next_level_cmd_payload_len;
  wire       [2:0]    iCache_1_next_level_cmd_payload_size;
  wire                sramBanks_2_sram_0_ports_rsp_valid;
  wire       [511:0]  sramBanks_2_sram_0_ports_rsp_payload_data;
  wire                sramBanks_2_sram_1_ports_rsp_valid;
  wire       [511:0]  sramBanks_2_sram_1_ports_rsp_payload_data;
  wire                sramBanks_2_sram_2_ports_rsp_valid;
  wire       [511:0]  sramBanks_2_sram_2_ports_rsp_payload_data;
  wire                sramBanks_2_sram_3_ports_rsp_valid;
  wire       [511:0]  sramBanks_2_sram_3_ports_rsp_payload_data;
  wire                dCache_1_stall;
  wire                dCache_1_cpu_cmd_ready;
  wire                dCache_1_cpu_rsp_valid;
  wire       [63:0]   dCache_1_cpu_rsp_payload_data;
  wire                dCache_1_sram_0_ports_cmd_valid;
  wire       [6:0]    dCache_1_sram_0_ports_cmd_payload_addr;
  wire       [7:0]    dCache_1_sram_0_ports_cmd_payload_wen;
  wire       [511:0]  dCache_1_sram_0_ports_cmd_payload_wdata;
  wire       [63:0]   dCache_1_sram_0_ports_cmd_payload_wstrb;
  wire                dCache_1_sram_1_ports_cmd_valid;
  wire       [6:0]    dCache_1_sram_1_ports_cmd_payload_addr;
  wire       [7:0]    dCache_1_sram_1_ports_cmd_payload_wen;
  wire       [511:0]  dCache_1_sram_1_ports_cmd_payload_wdata;
  wire       [63:0]   dCache_1_sram_1_ports_cmd_payload_wstrb;
  wire                dCache_1_sram_2_ports_cmd_valid;
  wire       [6:0]    dCache_1_sram_2_ports_cmd_payload_addr;
  wire       [7:0]    dCache_1_sram_2_ports_cmd_payload_wen;
  wire       [511:0]  dCache_1_sram_2_ports_cmd_payload_wdata;
  wire       [63:0]   dCache_1_sram_2_ports_cmd_payload_wstrb;
  wire                dCache_1_sram_3_ports_cmd_valid;
  wire       [6:0]    dCache_1_sram_3_ports_cmd_payload_addr;
  wire       [7:0]    dCache_1_sram_3_ports_cmd_payload_wen;
  wire       [511:0]  dCache_1_sram_3_ports_cmd_payload_wdata;
  wire       [63:0]   dCache_1_sram_3_ports_cmd_payload_wstrb;
  wire                dCache_1_next_level_cmd_valid;
  wire       [63:0]   dCache_1_next_level_cmd_payload_addr;
  wire       [3:0]    dCache_1_next_level_cmd_payload_len;
  wire       [2:0]    dCache_1_next_level_cmd_payload_size;
  wire                dCache_1_next_level_cmd_payload_wen;
  wire       [63:0]   dCache_1_next_level_cmd_payload_wdata;
  wire       [7:0]    dCache_1_next_level_cmd_payload_wstrb;
  wire                sramBanks_3_sram_0_ports_rsp_valid;
  wire       [511:0]  sramBanks_3_sram_0_ports_rsp_payload_data;
  wire                sramBanks_3_sram_1_ports_rsp_valid;
  wire       [511:0]  sramBanks_3_sram_1_ports_rsp_payload_data;
  wire                sramBanks_3_sram_2_ports_rsp_valid;
  wire       [511:0]  sramBanks_3_sram_2_ports_rsp_payload_data;
  wire                sramBanks_3_sram_3_ports_rsp_valid;
  wire       [511:0]  sramBanks_3_sram_3_ports_rsp_payload_data;
  wire       [11:0]   _zz__zz_decode_DecodePlugin_imm_2;
  wire       [11:0]   _zz__zz_decode_DecodePlugin_imm_4;
  wire       [19:0]   _zz__zz_decode_DecodePlugin_imm_6;
  wire       [31:0]   _zz__zz_decode_DecodePlugin_imm_8;
  wire       [63:0]   _zz_execute_ALUPlugin_add_result;
  wire       [63:0]   _zz_execute_ALUPlugin_add_result_1;
  wire       [63:0]   _zz_execute_ALUPlugin_sub_result;
  wire       [63:0]   _zz_execute_ALUPlugin_sub_result_1;
  wire       [63:0]   _zz_execute_ALUPlugin_slt_result;
  wire       [63:0]   _zz_execute_ALUPlugin_slt_result_1;
  wire       [63:0]   _zz_execute_ALUPlugin_sra_result;
  wire       [31:0]   _zz_execute_ALUPlugin_addw_result_2;
  wire       [31:0]   _zz_execute_ALUPlugin_subw_result_2;
  wire       [31:0]   _zz_execute_ALUPlugin_sraw_temp;
  wire       [63:0]   _zz_execute_ALUPlugin_blt_result;
  wire       [63:0]   _zz_execute_ALUPlugin_blt_result_1;
  wire       [63:0]   _zz_execute_ALUPlugin_bge_result;
  wire       [63:0]   _zz_execute_ALUPlugin_bge_result_1;
  wire       [63:0]   _zz_execute_ALUPlugin_pc_next;
  wire       [63:0]   _zz_execute_ALUPlugin_pc_next_1;
  wire       [63:0]   _zz_execute_ALUPlugin_pc_next_2;
  wire       [63:0]   _zz_execute_ALUPlugin_pc_next_3;
  wire       [63:0]   _zz_execute_ALUPlugin_pc_next_4;
  wire       [63:0]   _zz_execute_ALUPlugin_pc_next_5;
  wire       [63:0]   _zz_execute_ALUPlugin_pc_next_6;
  wire       [63:0]   _zz_execute_ALUPlugin_pc_next_7;
  wire       [63:0]   _zz_execute_ALUPlugin_pc_next_8;
  wire       [5:0]    _zz_memaccess_LSUPlugin_dcache_rdata;
  wire       [5:0]    _zz_memaccess_LSUPlugin_lsu_wdata;
  wire       [63:0]   writeback_RD;
  wire                memaccess_LSU_HOLD;
  wire                memaccess_TIMER_CEN;
  wire       [63:0]   memaccess_LSU_WDATA;
  wire                execute_INT_HOLD;
  wire       [63:0]   execute_REDIRECT_PC_NEXT;
  wire                execute_REDIRECT_VALID;
  wire                execute_IS_RET;
  wire                execute_IS_CALL;
  wire                execute_IS_JMP;
  wire       [6:0]    execute_BRANCH_HISTORY;
  wire                execute_BRANCH_TAKEN;
  wire                execute_BRANCH_OR_JUMP;
  wire                execute_BRANCH_OR_JALR;
  wire       [63:0]   execute_MEM_WDATA;
  wire       [63:0]   execute_ALU_RESULT;
  wire       [63:0]   decode_CSR_RDATA;
  wire                execute_CSR_WEN;
  wire                decode_CSR_WEN;
  wire       [11:0]   execute_CSR_ADDR;
  wire       [11:0]   decode_CSR_ADDR;
  wire       [3:0]    decode_CSR_CTRL;
  wire                execute_IS_STORE;
  wire                decode_IS_STORE;
  wire                execute_IS_LOAD;
  wire                decode_IS_LOAD;
  wire       [4:0]    writeback_RD_ADDR;
  wire       [4:0]    memaccess_RD_ADDR;
  wire       [4:0]    decode_RD_ADDR;
  wire                writeback_RD_WEN;
  wire                memaccess_RD_WEN;
  wire                execute_RD_WEN;
  wire                decode_RD_WEN;
  wire       [3:0]    execute_MEM_CTRL;
  wire       [3:0]    decode_MEM_CTRL;
  wire                decode_SRC2_IS_IMM;
  wire                decode_ALU_WORD;
  wire       [4:0]    decode_ALU_CTRL;
  wire       [4:0]    execute_RS2_ADDR;
  wire       [4:0]    decode_RS2_ADDR;
  wire       [4:0]    decode_RS1_ADDR;
  wire       [63:0]   decode_RS2;
  wire       [63:0]   decode_RS1;
  wire       [63:0]   decode_IMM;
  wire       [63:0]   fetch_INT_PC;
  wire                fetch_INT_EN;
  wire       [63:0]   fetch_PREDICT_PC;
  wire                decode_PREDICT_TAKEN;
  wire                fetch_PREDICT_TAKEN;
  wire                fetch_PREDICT_VALID;
  wire       [31:0]   memaccess_INSTRUCTION;
  wire       [31:0]   execute_INSTRUCTION;
  wire       [31:0]   fetch_INSTRUCTION;
  wire       [63:0]   decode_PC_NEXT;
  wire       [63:0]   fetch_PC_NEXT;
  wire       [63:0]   memaccess_PC;
  wire       [63:0]   fetch_PC;
  wire       [31:0]   writeback_INSTRUCTION;
  wire       [63:0]   writeback_PC;
  wire       [63:0]   writeback_ALU_RESULT;
  wire       [63:0]   writeback_LSU_RDATA;
  wire                writeback_IS_LOAD;
  wire       [3:0]    memaccess_MEM_CTRL;
  wire       [63:0]   memaccess_MEM_WDATA;
  wire                memaccess_IS_STORE;
  wire                memaccess_IS_LOAD;
  wire       [3:0]    execute_CSR_CTRL;
  wire       [63:0]   execute_SRC1;
  wire       [3:0]    _zz_ecall;
  wire       [11:0]   _zz_decode_to_execute_CSR_ADDR;
  wire                _zz_memaccess_arbitration_haltItself;
  wire                _zz_DecodePlugin_hazard_ctrl_rs1_from_mem;
  wire       [4:0]    _zz_DecodePlugin_hazard_rs2_from_mem;
  wire                _zz_DecodePlugin_hazard_rs1_from_mem;
  wire       [4:0]    _zz_DecodePlugin_hazard_rs1_from_mem_1;
  wire       [4:0]    _zz_DecodePlugin_hazard_rs1_from_mem_2;
  wire                _zz_DecodePlugin_hazard_rs1_from_mem_3;
  wire       [63:0]   execute_PC_NEXT;
  wire                execute_PREDICT_TAKEN;
  wire       [63:0]   execute_CSR_RDATA;
  wire                execute_ALU_WORD;
  wire                execute_CTRL_RS2_FROM_WB;
  wire                execute_CTRL_RS2_FROM_LOAD;
  wire                execute_CTRL_RS2_FROM_MEM;
  wire                execute_CTRL_RS1_FROM_WB;
  wire       [63:0]   _zz_execute_MEM_WDATA;
  wire                execute_CTRL_RS1_FROM_LOAD;
  wire       [63:0]   _zz_execute_MEM_WDATA_1;
  wire                execute_CTRL_RS1_FROM_MEM;
  wire       [63:0]   execute_RS2;
  wire                execute_RS2_FROM_WB;
  wire                execute_RS2_FROM_LOAD;
  wire                execute_RS2_FROM_MEM;
  wire       [63:0]   execute_IMM;
  wire                execute_SRC2_IS_IMM;
  wire       [63:0]   execute_RS1;
  wire                execute_RS1_FROM_WB;
  wire       [63:0]   memaccess_LSU_RDATA;
  wire                execute_RS1_FROM_LOAD;
  wire       [63:0]   memaccess_ALU_RESULT;
  wire                execute_RS1_FROM_MEM;
  wire       [63:0]   execute_PC;
  wire       [4:0]    execute_RS1_ADDR;
  wire       [4:0]    execute_RD_ADDR;
  wire       [4:0]    execute_ALU_CTRL;
  wire       [63:0]   _zz_execute_MEM_WDATA_2;
  wire       [4:0]    _zz_DecodePlugin_hazard_rs1_from_wb;
  wire                _zz_DecodePlugin_hazard_rs1_from_wb_1;
  wire       [31:0]   decode_INSTRUCTION;
  wire       [63:0]   decode_PC;
  wire       [63:0]   _zz_execute_to_memaccess_PC;
  wire       [63:0]   fetch_BPU_PC_NEXT;
  wire       [63:0]   _zz_pc_next;
  wire                when_FetchPlugin_l97;
  wire                fetch_BPU_BRANCH_TAKEN;
  wire                when_FetchPlugin_l94;
  wire                fetch_arbitration_haltItself;
  wire                fetch_arbitration_haltByOther;
  reg                 fetch_arbitration_removeIt;
  wire                fetch_arbitration_flushIt;
  wire                fetch_arbitration_flushNext;
  wire                fetch_arbitration_isValid;
  wire                fetch_arbitration_isStuck;
  wire                fetch_arbitration_isStuckByOthers;
  wire                fetch_arbitration_isFlushed;
  wire                fetch_arbitration_isMoving;
  wire                fetch_arbitration_isFiring;
  wire                decode_arbitration_haltItself;
  wire                decode_arbitration_haltByOther;
  reg                 decode_arbitration_removeIt;
  wire                decode_arbitration_flushIt;
  wire                decode_arbitration_flushNext;
  reg                 decode_arbitration_isValid;
  wire                decode_arbitration_isStuck;
  wire                decode_arbitration_isStuckByOthers;
  wire                decode_arbitration_isFlushed;
  wire                decode_arbitration_isMoving;
  wire                decode_arbitration_isFiring;
  wire                execute_arbitration_haltItself;
  wire                execute_arbitration_haltByOther;
  reg                 execute_arbitration_removeIt;
  wire                execute_arbitration_flushIt;
  wire                execute_arbitration_flushNext;
  reg                 execute_arbitration_isValid;
  wire                execute_arbitration_isStuck;
  wire                execute_arbitration_isStuckByOthers;
  wire                execute_arbitration_isFlushed;
  wire                execute_arbitration_isMoving;
  wire                execute_arbitration_isFiring;
  wire                memaccess_arbitration_haltItself;
  wire                memaccess_arbitration_haltByOther;
  reg                 memaccess_arbitration_removeIt;
  wire                memaccess_arbitration_flushIt;
  wire                memaccess_arbitration_flushNext;
  reg                 memaccess_arbitration_isValid;
  wire                memaccess_arbitration_isStuck;
  wire                memaccess_arbitration_isStuckByOthers;
  wire                memaccess_arbitration_isFlushed;
  wire                memaccess_arbitration_isMoving;
  wire                memaccess_arbitration_isFiring;
  wire                writeback_arbitration_haltItself;
  wire                writeback_arbitration_haltByOther;
  reg                 writeback_arbitration_removeIt;
  wire                writeback_arbitration_flushIt;
  wire                writeback_arbitration_flushNext;
  reg                 writeback_arbitration_isValid;
  wire                writeback_arbitration_isStuck;
  wire                writeback_arbitration_isStuckByOthers;
  wire                writeback_arbitration_isFlushed;
  wire                writeback_arbitration_isMoving;
  wire                writeback_arbitration_isFiring;
  wire                DecodePlugin_hazard_decode_rs1_req;
  wire                DecodePlugin_hazard_decode_rs2_req;
  wire       [4:0]    DecodePlugin_hazard_decode_rs1_addr;
  wire       [4:0]    DecodePlugin_hazard_decode_rs2_addr;
  wire                DecodePlugin_hazard_rs1_from_mem;
  wire                DecodePlugin_hazard_rs2_from_mem;
  wire                DecodePlugin_hazard_rs1_from_load;
  wire                DecodePlugin_hazard_rs2_from_load;
  wire                DecodePlugin_hazard_rs1_from_wb;
  wire                DecodePlugin_hazard_rs2_from_wb;
  wire                DecodePlugin_hazard_load_use;
  wire                DecodePlugin_hazard_ctrl_rs1_from_mem;
  wire                DecodePlugin_hazard_ctrl_rs2_from_mem;
  wire                DecodePlugin_hazard_ctrl_rs1_from_load;
  wire                DecodePlugin_hazard_ctrl_rs2_from_load;
  wire                DecodePlugin_hazard_ctrl_rs1_from_wb;
  wire                DecodePlugin_hazard_ctrl_rs2_from_wb;
  wire                DecodePlugin_hazard_ctrl_load_use;
  wire                ICachePlugin_icache_access_cmd_valid;
  wire                ICachePlugin_icache_access_cmd_ready;
  wire       [63:0]   ICachePlugin_icache_access_cmd_payload_addr;
  wire                ICachePlugin_icache_access_rsp_valid;
  wire       [31:0]   ICachePlugin_icache_access_rsp_payload_data;
  wire                DCachePlugin_dcache_access_cmd_valid;
  wire                DCachePlugin_dcache_access_cmd_ready;
  wire       [63:0]   DCachePlugin_dcache_access_cmd_payload_addr;
  wire                DCachePlugin_dcache_access_cmd_payload_wen;
  wire       [63:0]   DCachePlugin_dcache_access_cmd_payload_wdata;
  wire       [7:0]    DCachePlugin_dcache_access_cmd_payload_wstrb;
  wire                DCachePlugin_dcache_access_rsp_valid;
  wire       [63:0]   DCachePlugin_dcache_access_rsp_payload_data;
  wire                DCachePlugin_dcache_access_stall;
  reg        [63:0]   pc_next;
  reg                 fetch_valid;
  reg                 rsp_flush;
  wire                fetch_FetchPlugin_fetch_flush;
  wire                ICachePlugin_icache_access_cmd_fire;
  wire                fetch_FetchPlugin_bpu_predict_taken;
  wire                fetch_FetchPlugin_pc_in_stream_valid;
  wire                fetch_FetchPlugin_pc_in_stream_ready;
  wire       [63:0]   fetch_FetchPlugin_pc_in_stream_payload;
  wire                fetch_FetchPlugin_pc_out_stream_valid;
  wire                fetch_FetchPlugin_pc_out_stream_ready;
  wire       [63:0]   fetch_FetchPlugin_pc_out_stream_payload;
  wire                fetch_FetchPlugin_predict_taken_in_valid;
  wire                fetch_FetchPlugin_predict_taken_in_ready;
  wire                fetch_FetchPlugin_predict_taken_in_payload;
  wire                fetch_FetchPlugin_predict_taken_out_valid;
  wire                fetch_FetchPlugin_predict_taken_out_ready;
  wire                fetch_FetchPlugin_predict_taken_out_payload;
  wire                fetch_FetchPlugin_instruction_in_stream_valid;
  wire                fetch_FetchPlugin_instruction_in_stream_ready;
  wire       [31:0]   fetch_FetchPlugin_instruction_in_stream_payload;
  wire                fetch_FetchPlugin_instruction_out_stream_valid;
  wire                fetch_FetchPlugin_instruction_out_stream_ready;
  wire       [31:0]   fetch_FetchPlugin_instruction_out_stream_payload;
  wire                fetch_FetchPlugin_fifo_all_valid;
  wire       [1:0]    IDLE;
  wire       [1:0]    FETCH;
  wire       [1:0]    HALT;
  reg        [1:0]    fetch_state_next;
  reg        [1:0]    fetch_state;
  wire                when_FetchPlugin_l64;
  wire                ICachePlugin_icache_access_cmd_isStall;
  wire                when_FetchPlugin_l72;
  wire                when_FetchPlugin_l80;
  wire                when_FetchPlugin_l93;
  wire                when_FetchPlugin_l109;
  wire                ICachePlugin_icache_access_cmd_fire_1;
  wire                ICachePlugin_icache_access_cmd_fire_2;
  wire                ICachePlugin_icache_access_cmd_fire_3;
  wire                ICachePlugin_icache_access_cmd_fire_4;
  reg        [63:0]   decode_DecodePlugin_imm;
  wire       [63:0]   decode_DecodePlugin_rs1;
  wire       [63:0]   decode_DecodePlugin_rs2;
  wire                decode_DecodePlugin_rs1_req;
  wire                decode_DecodePlugin_rs2_req;
  wire       [4:0]    decode_DecodePlugin_rs1_addr;
  wire       [4:0]    decode_DecodePlugin_rs2_addr;
  wire                decode_DecodePlugin_rd_wen;
  wire       [4:0]    decode_DecodePlugin_rd_addr;
  reg        [4:0]    decode_DecodePlugin_alu_ctrl;
  wire                decode_DecodePlugin_alu_word;
  wire                decode_DecodePlugin_src2_is_imm;
  reg        [3:0]    decode_DecodePlugin_mem_ctrl;
  reg                 decode_DecodePlugin_is_load;
  reg                 decode_DecodePlugin_is_store;
  reg        [3:0]    decode_DecodePlugin_csr_ctrl;
  wire       [11:0]   decode_DecodePlugin_csr_addr;
  wire                decode_DecodePlugin_csr_wen;
  wire                when_DecodePlugin_l116;
  wire                _zz_decode_DecodePlugin_imm;
  reg        [51:0]   _zz_decode_DecodePlugin_imm_1;
  wire                _zz_decode_DecodePlugin_imm_2;
  reg        [51:0]   _zz_decode_DecodePlugin_imm_3;
  wire                _zz_decode_DecodePlugin_imm_4;
  reg        [50:0]   _zz_decode_DecodePlugin_imm_5;
  wire                _zz_decode_DecodePlugin_imm_6;
  reg        [42:0]   _zz_decode_DecodePlugin_imm_7;
  wire                _zz_decode_DecodePlugin_imm_8;
  reg        [31:0]   _zz_decode_DecodePlugin_imm_9;
  wire                _zz_decode_DecodePlugin_imm_10;
  reg        [51:0]   _zz_decode_DecodePlugin_imm_11;
  wire                when_DecodePlugin_l119;
  wire                when_DecodePlugin_l122;
  wire                when_DecodePlugin_l125;
  wire                when_DecodePlugin_l128;
  reg        [63:0]   execute_ALUPlugin_src1;
  reg        [63:0]   execute_ALUPlugin_src2;
  wire       [31:0]   execute_ALUPlugin_src1_word;
  wire       [31:0]   execute_ALUPlugin_src2_word;
  wire       [5:0]    execute_ALUPlugin_shift_bits;
  wire       [63:0]   execute_ALUPlugin_add_result;
  wire       [63:0]   execute_ALUPlugin_sub_result;
  wire                execute_ALUPlugin_slt_result;
  wire                execute_ALUPlugin_sltu_result;
  wire       [63:0]   execute_ALUPlugin_xor_result;
  wire       [63:0]   execute_ALUPlugin_sll_result;
  wire       [63:0]   execute_ALUPlugin_srl_result;
  wire       [63:0]   execute_ALUPlugin_sra_result;
  wire       [63:0]   execute_ALUPlugin_and_result;
  wire       [63:0]   execute_ALUPlugin_or_result;
  wire                _zz_execute_ALUPlugin_addw_result;
  reg        [31:0]   _zz_execute_ALUPlugin_addw_result_1;
  wire       [63:0]   execute_ALUPlugin_addw_result;
  wire                _zz_execute_ALUPlugin_subw_result;
  reg        [31:0]   _zz_execute_ALUPlugin_subw_result_1;
  wire       [63:0]   execute_ALUPlugin_subw_result;
  wire       [31:0]   execute_ALUPlugin_sllw_temp;
  wire                _zz_execute_ALUPlugin_sllw_result;
  reg        [31:0]   _zz_execute_ALUPlugin_sllw_result_1;
  wire       [63:0]   execute_ALUPlugin_sllw_result;
  wire       [31:0]   execute_ALUPlugin_srlw_temp;
  wire                _zz_execute_ALUPlugin_srlw_result;
  reg        [31:0]   _zz_execute_ALUPlugin_srlw_result_1;
  wire       [63:0]   execute_ALUPlugin_srlw_result;
  wire       [31:0]   execute_ALUPlugin_sraw_temp;
  wire                _zz_execute_ALUPlugin_sraw_result;
  reg        [31:0]   _zz_execute_ALUPlugin_sraw_result_1;
  wire       [63:0]   execute_ALUPlugin_sraw_result;
  reg        [63:0]   execute_ALUPlugin_alu_result;
  reg        [63:0]   execute_ALUPlugin_pc_next;
  wire                execute_ALUPlugin_jal;
  wire                execute_ALUPlugin_jalr;
  wire                execute_ALUPlugin_beq;
  wire                execute_ALUPlugin_bne;
  wire                execute_ALUPlugin_blt;
  wire                execute_ALUPlugin_bge;
  wire                execute_ALUPlugin_bltu;
  wire                execute_ALUPlugin_bgeu;
  wire                execute_ALUPlugin_branch_or_jalr;
  wire                execute_ALUPlugin_branch_or_jump;
  reg        [63:0]   execute_ALUPlugin_branch_src1;
  reg        [63:0]   execute_ALUPlugin_branch_src2;
  wire                execute_ALUPlugin_rd_is_link;
  wire                execute_ALUPlugin_rs1_is_link;
  reg                 execute_ALUPlugin_is_call;
  reg                 execute_ALUPlugin_is_ret;
  reg                 execute_ALUPlugin_is_jmp;
  reg        [63:0]   execute_ALUPlugin_redirect_pc_next;
  reg                 execute_ALUPlugin_redirect_valid;
  wire                when_AluPlugin_l77;
  wire                when_AluPlugin_l95;
  wire                when_AluPlugin_l146;
  wire                when_AluPlugin_l153;
  wire       [62:0]   _zz_execute_ALUPlugin_alu_result;
  wire       [62:0]   _zz_execute_ALUPlugin_alu_result_1;
  wire                when_AluPlugin_l169;
  wire                when_AluPlugin_l176;
  wire                when_AluPlugin_l183;
  wire                execute_ALUPlugin_beq_result;
  wire                execute_ALUPlugin_bne_result;
  wire                execute_ALUPlugin_blt_result;
  wire                execute_ALUPlugin_bge_result;
  wire                execute_ALUPlugin_bltu_result;
  wire                execute_ALUPlugin_bgeu_result;
  wire                execute_ALUPlugin_branch_taken;
  reg        [6:0]    execute_ALUPlugin_branch_history;
  wire                when_AluPlugin_l226;
  wire                when_AluPlugin_l234;
  wire                when_AluPlugin_l270;
  reg        [63:0]   execute_ExcepPlugin_csr_wdata;
  wire       [63:0]   execute_ExcepPlugin_csrrs_wdata;
  wire       [63:0]   execute_ExcepPlugin_csrrc_wdata;
  wire       [63:0]   execute_ExcepPlugin_csrrsi_wdata;
  wire       [63:0]   execute_ExcepPlugin_csrrci_wdata;
  wire       [63:0]   memaccess_LSUPlugin_cpu_addr;
  wire       [2:0]    memaccess_LSUPlugin_cpu_addr_offset;
  wire                memaccess_LSUPlugin_is_mem;
  wire                memaccess_LSUPlugin_is_timer;
  wire       [63:0]   memaccess_LSUPlugin_dcache_rdata;
  wire                _zz_memaccess_LSUPlugin_dcache_lb;
  reg        [55:0]   _zz_memaccess_LSUPlugin_dcache_lb_1;
  wire       [63:0]   memaccess_LSUPlugin_dcache_lb;
  reg        [55:0]   _zz_memaccess_LSUPlugin_dcache_lbu;
  wire       [63:0]   memaccess_LSUPlugin_dcache_lbu;
  wire                _zz_memaccess_LSUPlugin_dcache_lh;
  reg        [47:0]   _zz_memaccess_LSUPlugin_dcache_lh_1;
  wire       [63:0]   memaccess_LSUPlugin_dcache_lh;
  reg        [47:0]   _zz_memaccess_LSUPlugin_dcache_lhu;
  wire       [63:0]   memaccess_LSUPlugin_dcache_lhu;
  wire                _zz_memaccess_LSUPlugin_dcache_lw;
  reg        [31:0]   _zz_memaccess_LSUPlugin_dcache_lw_1;
  wire       [63:0]   memaccess_LSUPlugin_dcache_lw;
  reg        [31:0]   _zz_memaccess_LSUPlugin_dcache_lwu;
  wire       [63:0]   memaccess_LSUPlugin_dcache_lwu;
  reg        [63:0]   memaccess_LSUPlugin_dcache_data_load;
  wire                _zz_memaccess_LSUPlugin_dcache_sb;
  reg        [55:0]   _zz_memaccess_LSUPlugin_dcache_sb_1;
  wire       [63:0]   memaccess_LSUPlugin_dcache_sb;
  wire                _zz_memaccess_LSUPlugin_dcache_sh;
  reg        [47:0]   _zz_memaccess_LSUPlugin_dcache_sh_1;
  wire       [63:0]   memaccess_LSUPlugin_dcache_sh;
  wire                _zz_memaccess_LSUPlugin_dcache_sw;
  reg        [31:0]   _zz_memaccess_LSUPlugin_dcache_sw_1;
  wire       [63:0]   memaccess_LSUPlugin_dcache_sw;
  reg        [63:0]   memaccess_LSUPlugin_dcache_wdata;
  reg        [7:0]    memaccess_LSUPlugin_dcache_wstrb;
  wire                memaccess_LSUPlugin_lsu_ready;
  wire       [63:0]   memaccess_LSUPlugin_lsu_addr;
  wire       [63:0]   memaccess_LSUPlugin_lsu_rdata;
  wire       [63:0]   memaccess_LSUPlugin_lsu_wdata;
  wire                memaccess_LSUPlugin_lsu_wen;
  wire       [7:0]    memaccess_LSUPlugin_lsu_wstrb;
  reg        [7:0]    _zz_memaccess_LSUPlugin_dcache_wstrb;
  reg        [7:0]    _zz_memaccess_LSUPlugin_dcache_wstrb_1;
  reg        [7:0]    _zz_memaccess_LSUPlugin_dcache_wstrb_2;
  wire       [7:0]    _zz_memaccess_LSUPlugin_dcache_wstrb_3;
  reg                 _zz_when_DCachePlugin_l174;
  wire                when_DCachePlugin_l118;
  wire                dcache_ar_fire;
  wire                when_DCachePlugin_l141;
  wire                dcache_aw_fire;
  wire                when_DCachePlugin_l159;
  wire                dcache_w_fire;
  wire                when_DCachePlugin_l174;
  wire                dcache_aw_fire_1;
  wire                dcache_w_fire_1;
  wire                when_DCachePlugin_l175;
  wire                dcache_aw_fire_2;
  wire                dcache_w_fire_2;
  wire                when_DCachePlugin_l177;
  wire                dcache_aw_fire_3;
  wire                dcache_w_fire_3;
  wire                when_DCachePlugin_l182;
  wire                when_DCachePlugin_l181;
  wire                dcache_aw_fire_4;
  wire                dcache_w_fire_4;
  wire                dcache_aw_fire_5;
  wire                dcache_w_fire_5;
  wire                when_Pipeline_l127;
  reg        [63:0]   fetch_to_decode_PC;
  wire                when_Pipeline_l127_1;
  reg        [63:0]   decode_to_execute_PC;
  wire                when_Pipeline_l127_2;
  reg        [63:0]   execute_to_memaccess_PC;
  wire                when_Pipeline_l127_3;
  reg        [63:0]   memaccess_to_writeback_PC;
  wire                when_Pipeline_l127_4;
  reg        [63:0]   fetch_to_decode_PC_NEXT;
  wire                when_Pipeline_l127_5;
  reg        [63:0]   decode_to_execute_PC_NEXT;
  wire                when_Pipeline_l127_6;
  reg        [31:0]   fetch_to_decode_INSTRUCTION;
  wire                when_Pipeline_l127_7;
  reg        [31:0]   decode_to_execute_INSTRUCTION;
  wire                when_Pipeline_l127_8;
  reg        [31:0]   execute_to_memaccess_INSTRUCTION;
  wire                when_Pipeline_l127_9;
  reg        [31:0]   memaccess_to_writeback_INSTRUCTION;
  wire                when_Pipeline_l127_10;
  reg                 fetch_to_decode_PREDICT_TAKEN;
  wire                when_Pipeline_l127_11;
  reg                 decode_to_execute_PREDICT_TAKEN;
  wire                when_Pipeline_l127_12;
  reg        [63:0]   decode_to_execute_IMM;
  wire                when_Pipeline_l127_13;
  reg        [63:0]   decode_to_execute_RS1;
  wire                when_Pipeline_l127_14;
  reg        [63:0]   decode_to_execute_RS2;
  wire                when_Pipeline_l127_15;
  reg        [4:0]    decode_to_execute_RS1_ADDR;
  wire                when_Pipeline_l127_16;
  reg        [4:0]    decode_to_execute_RS2_ADDR;
  wire                when_Pipeline_l127_17;
  reg        [4:0]    decode_to_execute_ALU_CTRL;
  wire                when_Pipeline_l127_18;
  reg                 decode_to_execute_ALU_WORD;
  wire                when_Pipeline_l127_19;
  reg                 decode_to_execute_SRC2_IS_IMM;
  wire                when_Pipeline_l127_20;
  reg        [3:0]    decode_to_execute_MEM_CTRL;
  wire                when_Pipeline_l127_21;
  reg        [3:0]    execute_to_memaccess_MEM_CTRL;
  wire                when_Pipeline_l127_22;
  reg                 decode_to_execute_RD_WEN;
  wire                when_Pipeline_l127_23;
  reg                 execute_to_memaccess_RD_WEN;
  wire                when_Pipeline_l127_24;
  reg                 memaccess_to_writeback_RD_WEN;
  wire                when_Pipeline_l127_25;
  reg        [4:0]    decode_to_execute_RD_ADDR;
  wire                when_Pipeline_l127_26;
  reg        [4:0]    execute_to_memaccess_RD_ADDR;
  wire                when_Pipeline_l127_27;
  reg        [4:0]    memaccess_to_writeback_RD_ADDR;
  wire                when_Pipeline_l127_28;
  reg                 decode_to_execute_IS_LOAD;
  wire                when_Pipeline_l127_29;
  reg                 execute_to_memaccess_IS_LOAD;
  wire                when_Pipeline_l127_30;
  reg                 memaccess_to_writeback_IS_LOAD;
  wire                when_Pipeline_l127_31;
  reg                 decode_to_execute_IS_STORE;
  wire                when_Pipeline_l127_32;
  reg                 execute_to_memaccess_IS_STORE;
  wire                when_Pipeline_l127_33;
  reg        [3:0]    decode_to_execute_CSR_CTRL;
  wire                when_Pipeline_l127_34;
  reg        [11:0]   decode_to_execute_CSR_ADDR;
  wire                when_Pipeline_l127_35;
  reg                 decode_to_execute_CSR_WEN;
  wire                when_Pipeline_l127_36;
  reg        [63:0]   decode_to_execute_CSR_RDATA;
  wire                when_Pipeline_l127_37;
  reg        [63:0]   execute_to_memaccess_ALU_RESULT;
  wire                when_Pipeline_l127_38;
  reg        [63:0]   memaccess_to_writeback_ALU_RESULT;
  wire                when_Pipeline_l127_39;
  reg        [63:0]   execute_to_memaccess_MEM_WDATA;
  wire                when_Pipeline_l127_40;
  reg        [63:0]   memaccess_to_writeback_LSU_RDATA;
  wire                when_Pipeline_l163;
  wire                when_Pipeline_l166;
  wire                when_Pipeline_l163_1;
  wire                when_Pipeline_l166_1;
  wire                when_Pipeline_l163_2;
  wire                when_Pipeline_l166_2;
  wire                when_Pipeline_l163_3;
  wire                when_Pipeline_l166_3;
  function [55:0] zz__zz_memaccess_LSUPlugin_dcache_lbu(input dummy);
    begin
      zz__zz_memaccess_LSUPlugin_dcache_lbu[55] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[54] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[53] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[52] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[51] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[50] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[49] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[48] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[47] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[46] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[45] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[44] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[43] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[42] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[41] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[40] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[39] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[38] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[37] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[36] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[35] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[34] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[33] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[32] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[31] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[30] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[29] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[28] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[27] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[26] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[25] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[24] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[23] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[22] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[21] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[20] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[19] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[18] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[17] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[16] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[15] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[14] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[13] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[12] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[11] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[10] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[9] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[8] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[7] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[6] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[5] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[4] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[3] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[2] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[1] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lbu[0] = 1'b0;
    end
  endfunction
  wire [55:0] _zz_1;
  function [47:0] zz__zz_memaccess_LSUPlugin_dcache_lhu(input dummy);
    begin
      zz__zz_memaccess_LSUPlugin_dcache_lhu[47] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[46] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[45] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[44] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[43] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[42] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[41] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[40] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[39] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[38] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[37] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[36] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[35] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[34] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[33] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[32] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[31] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[30] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[29] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[28] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[27] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[26] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[25] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[24] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[23] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[22] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[21] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[20] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[19] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[18] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[17] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[16] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[15] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[14] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[13] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[12] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[11] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[10] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[9] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[8] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[7] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[6] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[5] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[4] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[3] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[2] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[1] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lhu[0] = 1'b0;
    end
  endfunction
  wire [47:0] _zz_2;
  function [31:0] zz__zz_memaccess_LSUPlugin_dcache_lwu(input dummy);
    begin
      zz__zz_memaccess_LSUPlugin_dcache_lwu[31] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[30] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[29] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[28] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[27] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[26] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[25] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[24] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[23] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[22] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[21] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[20] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[19] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[18] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[17] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[16] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[15] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[14] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[13] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[12] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[11] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[10] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[9] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[8] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[7] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[6] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[5] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[4] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[3] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[2] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[1] = 1'b0;
      zz__zz_memaccess_LSUPlugin_dcache_lwu[0] = 1'b0;
    end
  endfunction
  wire [31:0] _zz_3;
  function [7:0] zz__zz_memaccess_LSUPlugin_dcache_wstrb(input dummy);
    begin
      zz__zz_memaccess_LSUPlugin_dcache_wstrb = 8'h0;
      zz__zz_memaccess_LSUPlugin_dcache_wstrb[0] = 1'b1;
    end
  endfunction
  wire [7:0] _zz_4;
  function [7:0] zz__zz_memaccess_LSUPlugin_dcache_wstrb_1(input dummy);
    begin
      zz__zz_memaccess_LSUPlugin_dcache_wstrb_1 = 8'h0;
      zz__zz_memaccess_LSUPlugin_dcache_wstrb_1[1 : 0] = 2'b11;
    end
  endfunction
  wire [7:0] _zz_5;
  function [7:0] zz__zz_memaccess_LSUPlugin_dcache_wstrb_2(input dummy);
    begin
      zz__zz_memaccess_LSUPlugin_dcache_wstrb_2 = 8'h0;
      zz__zz_memaccess_LSUPlugin_dcache_wstrb_2[3 : 0] = 4'b1111;
    end
  endfunction
  wire [7:0] _zz_6;

  assign _zz__zz_decode_DecodePlugin_imm_2 = {decode_INSTRUCTION[31 : 25],decode_INSTRUCTION[11 : 7]};
  assign _zz__zz_decode_DecodePlugin_imm_4 = {{{decode_INSTRUCTION[31],decode_INSTRUCTION[7]},decode_INSTRUCTION[30 : 25]},decode_INSTRUCTION[11 : 8]};
  assign _zz__zz_decode_DecodePlugin_imm_6 = {{{decode_INSTRUCTION[31],decode_INSTRUCTION[19 : 12]},decode_INSTRUCTION[20]},decode_INSTRUCTION[30 : 21]};
  assign _zz__zz_decode_DecodePlugin_imm_8 = {decode_INSTRUCTION[31 : 12],12'h0};
  assign _zz_execute_ALUPlugin_add_result = execute_ALUPlugin_src1;
  assign _zz_execute_ALUPlugin_add_result_1 = execute_ALUPlugin_src2;
  assign _zz_execute_ALUPlugin_sub_result = execute_ALUPlugin_src1;
  assign _zz_execute_ALUPlugin_sub_result_1 = execute_ALUPlugin_src2;
  assign _zz_execute_ALUPlugin_slt_result = execute_ALUPlugin_src1;
  assign _zz_execute_ALUPlugin_slt_result_1 = execute_ALUPlugin_src2;
  assign _zz_execute_ALUPlugin_sra_result = execute_ALUPlugin_src1;
  assign _zz_execute_ALUPlugin_addw_result_2 = execute_ALUPlugin_add_result[31 : 0];
  assign _zz_execute_ALUPlugin_subw_result_2 = execute_ALUPlugin_sub_result[31 : 0];
  assign _zz_execute_ALUPlugin_sraw_temp = execute_ALUPlugin_src1_word;
  assign _zz_execute_ALUPlugin_blt_result = execute_ALUPlugin_branch_src1;
  assign _zz_execute_ALUPlugin_blt_result_1 = execute_ALUPlugin_branch_src2;
  assign _zz_execute_ALUPlugin_bge_result = execute_ALUPlugin_branch_src2;
  assign _zz_execute_ALUPlugin_bge_result_1 = execute_ALUPlugin_branch_src1;
  assign _zz_execute_ALUPlugin_pc_next = (_zz_execute_ALUPlugin_pc_next_1 & _zz_execute_ALUPlugin_pc_next_4);
  assign _zz_execute_ALUPlugin_pc_next_1 = ($signed(_zz_execute_ALUPlugin_pc_next_2) + $signed(_zz_execute_ALUPlugin_pc_next_3));
  assign _zz_execute_ALUPlugin_pc_next_2 = execute_ALUPlugin_branch_src1;
  assign _zz_execute_ALUPlugin_pc_next_3 = execute_IMM;
  assign _zz_execute_ALUPlugin_pc_next_4 = (~ _zz_execute_ALUPlugin_pc_next_5);
  assign _zz_execute_ALUPlugin_pc_next_5 = 64'h0000000000000001;
  assign _zz_execute_ALUPlugin_pc_next_6 = ($signed(_zz_execute_ALUPlugin_pc_next_7) + $signed(_zz_execute_ALUPlugin_pc_next_8));
  assign _zz_execute_ALUPlugin_pc_next_7 = execute_PC;
  assign _zz_execute_ALUPlugin_pc_next_8 = execute_IMM;
  assign _zz_memaccess_LSUPlugin_dcache_rdata = ({3'd0,memaccess_LSUPlugin_cpu_addr_offset} <<< 3);
  assign _zz_memaccess_LSUPlugin_lsu_wdata = ({3'd0,memaccess_LSUPlugin_cpu_addr_offset} <<< 3);
  FIFO fetch_FetchPlugin_pc_stream_fifo (
    .ports_s_ports_valid   (fetch_FetchPlugin_pc_in_stream_valid                        ), //i
    .ports_s_ports_ready   (fetch_FetchPlugin_pc_stream_fifo_ports_s_ports_ready        ), //o
    .ports_s_ports_payload (fetch_FetchPlugin_pc_in_stream_payload[63:0]                ), //i
    .ports_m_ports_valid   (fetch_FetchPlugin_pc_stream_fifo_ports_m_ports_valid        ), //o
    .ports_m_ports_ready   (fetch_FetchPlugin_pc_out_stream_ready                       ), //i
    .ports_m_ports_payload (fetch_FetchPlugin_pc_stream_fifo_ports_m_ports_payload[63:0]), //o
    .flush                 (fetch_FetchPlugin_fetch_flush                               ), //i
    .next_payload          (fetch_FetchPlugin_pc_stream_fifo_next_payload[63:0]         ), //o
    .next_valid            (fetch_FetchPlugin_pc_stream_fifo_next_valid                 ), //o
    .clk                   (clk                                                         ), //i
    .reset                 (reset                                                       )  //i
  );
  FIFO_1 fetch_FetchPlugin_predict_taken_fifo (
    .ports_s_ports_valid   (fetch_FetchPlugin_predict_taken_in_valid                  ), //i
    .ports_s_ports_ready   (fetch_FetchPlugin_predict_taken_fifo_ports_s_ports_ready  ), //o
    .ports_s_ports_payload (fetch_FetchPlugin_predict_taken_in_payload                ), //i
    .ports_m_ports_valid   (fetch_FetchPlugin_predict_taken_fifo_ports_m_ports_valid  ), //o
    .ports_m_ports_ready   (fetch_FetchPlugin_predict_taken_out_ready                 ), //i
    .ports_m_ports_payload (fetch_FetchPlugin_predict_taken_fifo_ports_m_ports_payload), //o
    .flush                 (fetch_FetchPlugin_fetch_flush                             ), //i
    .clk                   (clk                                                       ), //i
    .reset                 (reset                                                     )  //i
  );
  FIFO_2 fetch_FetchPlugin_instruction_stream_fifo (
    .ports_s_ports_valid   (fetch_FetchPlugin_instruction_in_stream_valid                        ), //i
    .ports_s_ports_ready   (fetch_FetchPlugin_instruction_stream_fifo_ports_s_ports_ready        ), //o
    .ports_s_ports_payload (fetch_FetchPlugin_instruction_in_stream_payload[31:0]                ), //i
    .ports_m_ports_valid   (fetch_FetchPlugin_instruction_stream_fifo_ports_m_ports_valid        ), //o
    .ports_m_ports_ready   (fetch_FetchPlugin_instruction_out_stream_ready                       ), //i
    .ports_m_ports_payload (fetch_FetchPlugin_instruction_stream_fifo_ports_m_ports_payload[31:0]), //o
    .flush                 (fetch_FetchPlugin_fetch_flush                                        ), //i
    .clk                   (clk                                                                  ), //i
    .reset                 (reset                                                                )  //i
  );
  gshare_predictor gshare_predictor_1 (
    .predict_pc         (fetch_PREDICT_PC[63:0]                  ), //i
    .predict_valid      (fetch_PREDICT_VALID                     ), //i
    .predict_taken      (gshare_predictor_1_predict_taken        ), //o
    .predict_history    (gshare_predictor_1_predict_history[6:0] ), //o
    .predict_pc_next    (gshare_predictor_1_predict_pc_next[63:0]), //o
    .train_valid        (execute_BRANCH_OR_JUMP                  ), //i
    .train_taken        (execute_BRANCH_TAKEN                    ), //i
    .train_mispredicted (when_FetchPlugin_l97                    ), //i
    .train_history      (execute_BRANCH_HISTORY[6:0]             ), //i
    .train_pc           (_zz_execute_to_memaccess_PC[63:0]       ), //i
    .train_pc_next      (_zz_pc_next[63:0]                       ), //i
    .train_is_call      (execute_IS_CALL                         ), //i
    .train_is_ret       (execute_IS_RET                          ), //i
    .train_is_jmp       (execute_IS_JMP                          ), //i
    .clk                (clk                                     ), //i
    .reset              (reset                                   )  //i
  );
  RegFileModule regFileModule_1 (
    .read_ports_rs1_value (regFileModule_1_read_ports_rs1_value[63:0]), //o
    .read_ports_rs2_value (regFileModule_1_read_ports_rs2_value[63:0]), //o
    .read_ports_rs1_addr  (decode_DecodePlugin_rs1_addr[4:0]         ), //i
    .read_ports_rs2_addr  (decode_DecodePlugin_rs2_addr[4:0]         ), //i
    .read_ports_rs1_req   (decode_DecodePlugin_rs1_req               ), //i
    .read_ports_rs2_req   (decode_DecodePlugin_rs2_req               ), //i
    .write_ports_rd_value (_zz_execute_MEM_WDATA_2[63:0]             ), //i
    .write_ports_rd_addr  (_zz_DecodePlugin_hazard_rs1_from_wb[4:0]  ), //i
    .write_ports_rd_wen   (regFileModule_1_write_ports_rd_wen        ), //i
    .clk                  (clk                                       ), //i
    .reset                (reset                                     )  //i
  );
  CsrRegfile csrRegfile_1 (
    .cpu_ports_waddr            (execute_CSR_ADDR[11:0]                 ), //i
    .cpu_ports_wen              (execute_CSR_WEN                        ), //i
    .cpu_ports_wdata            (execute_ExcepPlugin_csr_wdata[63:0]    ), //i
    .cpu_ports_raddr            (_zz_decode_to_execute_CSR_ADDR[11:0]   ), //i
    .cpu_ports_rdata            (csrRegfile_1_cpu_ports_rdata[63:0]     ), //o
    .clint_ports_mepc_wen       (clint_1_csr_ports_mepc_wen             ), //i
    .clint_ports_mepc_wdata     (clint_1_csr_ports_mepc_wdata[63:0]     ), //i
    .clint_ports_mcause_wen     (clint_1_csr_ports_mcause_wen           ), //i
    .clint_ports_mcause_wdata   (clint_1_csr_ports_mcause_wdata[63:0]   ), //i
    .clint_ports_mstatus_wen    (clint_1_csr_ports_mstatus_wen          ), //i
    .clint_ports_mstatus_wdata  (clint_1_csr_ports_mstatus_wdata[63:0]  ), //i
    .clint_ports_mtvec          (csrRegfile_1_clint_ports_mtvec[63:0]   ), //o
    .clint_ports_mepc           (csrRegfile_1_clint_ports_mepc[63:0]    ), //o
    .clint_ports_mstatus        (csrRegfile_1_clint_ports_mstatus[63:0] ), //o
    .clint_ports_global_int_en  (csrRegfile_1_clint_ports_global_int_en ), //o
    .clint_ports_mtime_int_en   (csrRegfile_1_clint_ports_mtime_int_en  ), //o
    .clint_ports_mtime_int_pend (csrRegfile_1_clint_ports_mtime_int_pend), //o
    .timer_int                  (timer_1_timer_int                      ), //i
    .clk                        (clk                                    ), //i
    .reset                      (reset                                  )  //i
  );
  Clint clint_1 (
    .pc                       (_zz_execute_to_memaccess_PC[63:0]      ), //i
    .pc_next                  (_zz_pc_next[63:0]                      ), //i
    .pc_next_valid            (when_FetchPlugin_l97                   ), //i
    .instruction_valid        (execute_arbitration_isValid            ), //i
    .csr_ports_mepc_wen       (clint_1_csr_ports_mepc_wen             ), //o
    .csr_ports_mepc_wdata     (clint_1_csr_ports_mepc_wdata[63:0]     ), //o
    .csr_ports_mcause_wen     (clint_1_csr_ports_mcause_wen           ), //o
    .csr_ports_mcause_wdata   (clint_1_csr_ports_mcause_wdata[63:0]   ), //o
    .csr_ports_mstatus_wen    (clint_1_csr_ports_mstatus_wen          ), //o
    .csr_ports_mstatus_wdata  (clint_1_csr_ports_mstatus_wdata[63:0]  ), //o
    .csr_ports_mtvec          (csrRegfile_1_clint_ports_mtvec[63:0]   ), //i
    .csr_ports_mepc           (csrRegfile_1_clint_ports_mepc[63:0]    ), //i
    .csr_ports_mstatus        (csrRegfile_1_clint_ports_mstatus[63:0] ), //i
    .csr_ports_global_int_en  (csrRegfile_1_clint_ports_global_int_en ), //i
    .csr_ports_mtime_int_en   (csrRegfile_1_clint_ports_mtime_int_en  ), //i
    .csr_ports_mtime_int_pend (csrRegfile_1_clint_ports_mtime_int_pend), //i
    .timer_int                (timer_1_timer_int                      ), //i
    .int_en                   (clint_1_int_en                         ), //o
    .int_pc                   (clint_1_int_pc[63:0]                   ), //o
    .int_hold                 (clint_1_int_hold                       ), //o
    .ecall                    (clint_1_ecall                          ), //i
    .ebreak                   (clint_1_ebreak                         ), //i
    .mret                     (clint_1_mret                           ), //i
    .clk                      (clk                                    ), //i
    .reset                    (reset                                  )  //i
  );
  Timer timer_1 (
    .cen       (memaccess_TIMER_CEN      ), //i
    .wen       (memaccess_IS_STORE       ), //i
    .addr      (timer_1_addr[63:0]       ), //i
    .wdata     (memaccess_LSU_WDATA[63:0]), //i
    .rdata     (timer_1_rdata[63:0]      ), //o
    .timer_int (timer_1_timer_int        ), //o
    .clk       (clk                      ), //i
    .reset     (reset                    )  //i
  );
  ICache iCache_1 (
    .flush                           (1'b0                                             ), //i
    .cpu_cmd_valid                   (ICachePlugin_icache_access_cmd_valid             ), //i
    .cpu_cmd_ready                   (iCache_1_cpu_cmd_ready                           ), //o
    .cpu_cmd_payload_addr            (ICachePlugin_icache_access_cmd_payload_addr[63:0]), //i
    .cpu_rsp_valid                   (iCache_1_cpu_rsp_valid                           ), //o
    .cpu_rsp_payload_data            (iCache_1_cpu_rsp_payload_data[31:0]              ), //o
    .sram_0_ports_cmd_valid          (iCache_1_sram_0_ports_cmd_valid                  ), //o
    .sram_0_ports_cmd_payload_addr   (iCache_1_sram_0_ports_cmd_payload_addr[6:0]      ), //o
    .sram_0_ports_cmd_payload_wen    (iCache_1_sram_0_ports_cmd_payload_wen[15:0]      ), //o
    .sram_0_ports_cmd_payload_wdata  (iCache_1_sram_0_ports_cmd_payload_wdata[511:0]   ), //o
    .sram_0_ports_cmd_payload_wstrb  (iCache_1_sram_0_ports_cmd_payload_wstrb[63:0]    ), //o
    .sram_0_ports_rsp_valid          (sramBanks_2_sram_0_ports_rsp_valid               ), //i
    .sram_0_ports_rsp_payload_data   (sramBanks_2_sram_0_ports_rsp_payload_data[511:0] ), //i
    .sram_1_ports_cmd_valid          (iCache_1_sram_1_ports_cmd_valid                  ), //o
    .sram_1_ports_cmd_payload_addr   (iCache_1_sram_1_ports_cmd_payload_addr[6:0]      ), //o
    .sram_1_ports_cmd_payload_wen    (iCache_1_sram_1_ports_cmd_payload_wen[15:0]      ), //o
    .sram_1_ports_cmd_payload_wdata  (iCache_1_sram_1_ports_cmd_payload_wdata[511:0]   ), //o
    .sram_1_ports_cmd_payload_wstrb  (iCache_1_sram_1_ports_cmd_payload_wstrb[63:0]    ), //o
    .sram_1_ports_rsp_valid          (sramBanks_2_sram_1_ports_rsp_valid               ), //i
    .sram_1_ports_rsp_payload_data   (sramBanks_2_sram_1_ports_rsp_payload_data[511:0] ), //i
    .sram_2_ports_cmd_valid          (iCache_1_sram_2_ports_cmd_valid                  ), //o
    .sram_2_ports_cmd_payload_addr   (iCache_1_sram_2_ports_cmd_payload_addr[6:0]      ), //o
    .sram_2_ports_cmd_payload_wen    (iCache_1_sram_2_ports_cmd_payload_wen[15:0]      ), //o
    .sram_2_ports_cmd_payload_wdata  (iCache_1_sram_2_ports_cmd_payload_wdata[511:0]   ), //o
    .sram_2_ports_cmd_payload_wstrb  (iCache_1_sram_2_ports_cmd_payload_wstrb[63:0]    ), //o
    .sram_2_ports_rsp_valid          (sramBanks_2_sram_2_ports_rsp_valid               ), //i
    .sram_2_ports_rsp_payload_data   (sramBanks_2_sram_2_ports_rsp_payload_data[511:0] ), //i
    .sram_3_ports_cmd_valid          (iCache_1_sram_3_ports_cmd_valid                  ), //o
    .sram_3_ports_cmd_payload_addr   (iCache_1_sram_3_ports_cmd_payload_addr[6:0]      ), //o
    .sram_3_ports_cmd_payload_wen    (iCache_1_sram_3_ports_cmd_payload_wen[15:0]      ), //o
    .sram_3_ports_cmd_payload_wdata  (iCache_1_sram_3_ports_cmd_payload_wdata[511:0]   ), //o
    .sram_3_ports_cmd_payload_wstrb  (iCache_1_sram_3_ports_cmd_payload_wstrb[63:0]    ), //o
    .sram_3_ports_rsp_valid          (sramBanks_2_sram_3_ports_rsp_valid               ), //i
    .sram_3_ports_rsp_payload_data   (sramBanks_2_sram_3_ports_rsp_payload_data[511:0] ), //i
    .sram_4_ports_cmd_valid          (iCache_1_sram_4_ports_cmd_valid                  ), //o
    .sram_4_ports_cmd_payload_addr   (iCache_1_sram_4_ports_cmd_payload_addr[6:0]      ), //o
    .sram_4_ports_cmd_payload_wen    (iCache_1_sram_4_ports_cmd_payload_wen[15:0]      ), //o
    .sram_4_ports_cmd_payload_wdata  (iCache_1_sram_4_ports_cmd_payload_wdata[511:0]   ), //o
    .sram_4_ports_cmd_payload_wstrb  (iCache_1_sram_4_ports_cmd_payload_wstrb[63:0]    ), //o
    .sram_4_ports_rsp_valid          (iCache_1_sram_4_ports_rsp_valid                  ), //i
    .sram_4_ports_rsp_payload_data   (iCache_1_sram_4_ports_rsp_payload_data[511:0]    ), //i
    .sram_5_ports_cmd_valid          (iCache_1_sram_5_ports_cmd_valid                  ), //o
    .sram_5_ports_cmd_payload_addr   (iCache_1_sram_5_ports_cmd_payload_addr[6:0]      ), //o
    .sram_5_ports_cmd_payload_wen    (iCache_1_sram_5_ports_cmd_payload_wen[15:0]      ), //o
    .sram_5_ports_cmd_payload_wdata  (iCache_1_sram_5_ports_cmd_payload_wdata[511:0]   ), //o
    .sram_5_ports_cmd_payload_wstrb  (iCache_1_sram_5_ports_cmd_payload_wstrb[63:0]    ), //o
    .sram_5_ports_rsp_valid          (iCache_1_sram_5_ports_rsp_valid                  ), //i
    .sram_5_ports_rsp_payload_data   (iCache_1_sram_5_ports_rsp_payload_data[511:0]    ), //i
    .sram_6_ports_cmd_valid          (iCache_1_sram_6_ports_cmd_valid                  ), //o
    .sram_6_ports_cmd_payload_addr   (iCache_1_sram_6_ports_cmd_payload_addr[6:0]      ), //o
    .sram_6_ports_cmd_payload_wen    (iCache_1_sram_6_ports_cmd_payload_wen[15:0]      ), //o
    .sram_6_ports_cmd_payload_wdata  (iCache_1_sram_6_ports_cmd_payload_wdata[511:0]   ), //o
    .sram_6_ports_cmd_payload_wstrb  (iCache_1_sram_6_ports_cmd_payload_wstrb[63:0]    ), //o
    .sram_6_ports_rsp_valid          (iCache_1_sram_6_ports_rsp_valid                  ), //i
    .sram_6_ports_rsp_payload_data   (iCache_1_sram_6_ports_rsp_payload_data[511:0]    ), //i
    .sram_7_ports_cmd_valid          (iCache_1_sram_7_ports_cmd_valid                  ), //o
    .sram_7_ports_cmd_payload_addr   (iCache_1_sram_7_ports_cmd_payload_addr[6:0]      ), //o
    .sram_7_ports_cmd_payload_wen    (iCache_1_sram_7_ports_cmd_payload_wen[15:0]      ), //o
    .sram_7_ports_cmd_payload_wdata  (iCache_1_sram_7_ports_cmd_payload_wdata[511:0]   ), //o
    .sram_7_ports_cmd_payload_wstrb  (iCache_1_sram_7_ports_cmd_payload_wstrb[63:0]    ), //o
    .sram_7_ports_rsp_valid          (iCache_1_sram_7_ports_rsp_valid                  ), //i
    .sram_7_ports_rsp_payload_data   (iCache_1_sram_7_ports_rsp_payload_data[511:0]    ), //i
    .sram_8_ports_cmd_valid          (iCache_1_sram_8_ports_cmd_valid                  ), //o
    .sram_8_ports_cmd_payload_addr   (iCache_1_sram_8_ports_cmd_payload_addr[6:0]      ), //o
    .sram_8_ports_cmd_payload_wen    (iCache_1_sram_8_ports_cmd_payload_wen[15:0]      ), //o
    .sram_8_ports_cmd_payload_wdata  (iCache_1_sram_8_ports_cmd_payload_wdata[511:0]   ), //o
    .sram_8_ports_cmd_payload_wstrb  (iCache_1_sram_8_ports_cmd_payload_wstrb[63:0]    ), //o
    .sram_8_ports_rsp_valid          (iCache_1_sram_8_ports_rsp_valid                  ), //i
    .sram_8_ports_rsp_payload_data   (iCache_1_sram_8_ports_rsp_payload_data[511:0]    ), //i
    .sram_9_ports_cmd_valid          (iCache_1_sram_9_ports_cmd_valid                  ), //o
    .sram_9_ports_cmd_payload_addr   (iCache_1_sram_9_ports_cmd_payload_addr[6:0]      ), //o
    .sram_9_ports_cmd_payload_wen    (iCache_1_sram_9_ports_cmd_payload_wen[15:0]      ), //o
    .sram_9_ports_cmd_payload_wdata  (iCache_1_sram_9_ports_cmd_payload_wdata[511:0]   ), //o
    .sram_9_ports_cmd_payload_wstrb  (iCache_1_sram_9_ports_cmd_payload_wstrb[63:0]    ), //o
    .sram_9_ports_rsp_valid          (iCache_1_sram_9_ports_rsp_valid                  ), //i
    .sram_9_ports_rsp_payload_data   (iCache_1_sram_9_ports_rsp_payload_data[511:0]    ), //i
    .sram_10_ports_cmd_valid         (iCache_1_sram_10_ports_cmd_valid                 ), //o
    .sram_10_ports_cmd_payload_addr  (iCache_1_sram_10_ports_cmd_payload_addr[6:0]     ), //o
    .sram_10_ports_cmd_payload_wen   (iCache_1_sram_10_ports_cmd_payload_wen[15:0]     ), //o
    .sram_10_ports_cmd_payload_wdata (iCache_1_sram_10_ports_cmd_payload_wdata[511:0]  ), //o
    .sram_10_ports_cmd_payload_wstrb (iCache_1_sram_10_ports_cmd_payload_wstrb[63:0]   ), //o
    .sram_10_ports_rsp_valid         (iCache_1_sram_10_ports_rsp_valid                 ), //i
    .sram_10_ports_rsp_payload_data  (iCache_1_sram_10_ports_rsp_payload_data[511:0]   ), //i
    .sram_11_ports_cmd_valid         (iCache_1_sram_11_ports_cmd_valid                 ), //o
    .sram_11_ports_cmd_payload_addr  (iCache_1_sram_11_ports_cmd_payload_addr[6:0]     ), //o
    .sram_11_ports_cmd_payload_wen   (iCache_1_sram_11_ports_cmd_payload_wen[15:0]     ), //o
    .sram_11_ports_cmd_payload_wdata (iCache_1_sram_11_ports_cmd_payload_wdata[511:0]  ), //o
    .sram_11_ports_cmd_payload_wstrb (iCache_1_sram_11_ports_cmd_payload_wstrb[63:0]   ), //o
    .sram_11_ports_rsp_valid         (iCache_1_sram_11_ports_rsp_valid                 ), //i
    .sram_11_ports_rsp_payload_data  (iCache_1_sram_11_ports_rsp_payload_data[511:0]   ), //i
    .sram_12_ports_cmd_valid         (iCache_1_sram_12_ports_cmd_valid                 ), //o
    .sram_12_ports_cmd_payload_addr  (iCache_1_sram_12_ports_cmd_payload_addr[6:0]     ), //o
    .sram_12_ports_cmd_payload_wen   (iCache_1_sram_12_ports_cmd_payload_wen[15:0]     ), //o
    .sram_12_ports_cmd_payload_wdata (iCache_1_sram_12_ports_cmd_payload_wdata[511:0]  ), //o
    .sram_12_ports_cmd_payload_wstrb (iCache_1_sram_12_ports_cmd_payload_wstrb[63:0]   ), //o
    .sram_12_ports_rsp_valid         (iCache_1_sram_12_ports_rsp_valid                 ), //i
    .sram_12_ports_rsp_payload_data  (iCache_1_sram_12_ports_rsp_payload_data[511:0]   ), //i
    .sram_13_ports_cmd_valid         (iCache_1_sram_13_ports_cmd_valid                 ), //o
    .sram_13_ports_cmd_payload_addr  (iCache_1_sram_13_ports_cmd_payload_addr[6:0]     ), //o
    .sram_13_ports_cmd_payload_wen   (iCache_1_sram_13_ports_cmd_payload_wen[15:0]     ), //o
    .sram_13_ports_cmd_payload_wdata (iCache_1_sram_13_ports_cmd_payload_wdata[511:0]  ), //o
    .sram_13_ports_cmd_payload_wstrb (iCache_1_sram_13_ports_cmd_payload_wstrb[63:0]   ), //o
    .sram_13_ports_rsp_valid         (iCache_1_sram_13_ports_rsp_valid                 ), //i
    .sram_13_ports_rsp_payload_data  (iCache_1_sram_13_ports_rsp_payload_data[511:0]   ), //i
    .sram_14_ports_cmd_valid         (iCache_1_sram_14_ports_cmd_valid                 ), //o
    .sram_14_ports_cmd_payload_addr  (iCache_1_sram_14_ports_cmd_payload_addr[6:0]     ), //o
    .sram_14_ports_cmd_payload_wen   (iCache_1_sram_14_ports_cmd_payload_wen[15:0]     ), //o
    .sram_14_ports_cmd_payload_wdata (iCache_1_sram_14_ports_cmd_payload_wdata[511:0]  ), //o
    .sram_14_ports_cmd_payload_wstrb (iCache_1_sram_14_ports_cmd_payload_wstrb[63:0]   ), //o
    .sram_14_ports_rsp_valid         (iCache_1_sram_14_ports_rsp_valid                 ), //i
    .sram_14_ports_rsp_payload_data  (iCache_1_sram_14_ports_rsp_payload_data[511:0]   ), //i
    .sram_15_ports_cmd_valid         (iCache_1_sram_15_ports_cmd_valid                 ), //o
    .sram_15_ports_cmd_payload_addr  (iCache_1_sram_15_ports_cmd_payload_addr[6:0]     ), //o
    .sram_15_ports_cmd_payload_wen   (iCache_1_sram_15_ports_cmd_payload_wen[15:0]     ), //o
    .sram_15_ports_cmd_payload_wdata (iCache_1_sram_15_ports_cmd_payload_wdata[511:0]  ), //o
    .sram_15_ports_cmd_payload_wstrb (iCache_1_sram_15_ports_cmd_payload_wstrb[63:0]   ), //o
    .sram_15_ports_rsp_valid         (iCache_1_sram_15_ports_rsp_valid                 ), //i
    .sram_15_ports_rsp_payload_data  (iCache_1_sram_15_ports_rsp_payload_data[511:0]   ), //i
    .next_level_cmd_valid            (iCache_1_next_level_cmd_valid                    ), //o
    .next_level_cmd_ready            (icache_ar_ready                                  ), //i
    .next_level_cmd_payload_addr     (iCache_1_next_level_cmd_payload_addr[63:0]       ), //o
    .next_level_cmd_payload_len      (iCache_1_next_level_cmd_payload_len[3:0]         ), //o
    .next_level_cmd_payload_size     (iCache_1_next_level_cmd_payload_size[2:0]        ), //o
    .next_level_rsp_valid            (icache_r_valid                                   ), //i
    .next_level_rsp_payload_data     (icache_r_payload_data[63:0]                      ), //i
    .clk                             (clk                                              ), //i
    .reset                           (reset                                            )  //i
  );
  SramBanks sramBanks_2 (
    .sram_0_ports_cmd_valid         (iCache_1_sram_0_ports_cmd_valid                 ), //i
    .sram_0_ports_cmd_payload_addr  (iCache_1_sram_0_ports_cmd_payload_addr[6:0]     ), //i
    .sram_0_ports_cmd_payload_wen   (iCache_1_sram_0_ports_cmd_payload_wen[15:0]     ), //i
    .sram_0_ports_cmd_payload_wdata (iCache_1_sram_0_ports_cmd_payload_wdata[511:0]  ), //i
    .sram_0_ports_cmd_payload_wstrb (iCache_1_sram_0_ports_cmd_payload_wstrb[63:0]   ), //i
    .sram_0_ports_rsp_valid         (sramBanks_2_sram_0_ports_rsp_valid              ), //o
    .sram_0_ports_rsp_payload_data  (sramBanks_2_sram_0_ports_rsp_payload_data[511:0]), //o
    .sram_1_ports_cmd_valid         (iCache_1_sram_1_ports_cmd_valid                 ), //i
    .sram_1_ports_cmd_payload_addr  (iCache_1_sram_1_ports_cmd_payload_addr[6:0]     ), //i
    .sram_1_ports_cmd_payload_wen   (iCache_1_sram_1_ports_cmd_payload_wen[15:0]     ), //i
    .sram_1_ports_cmd_payload_wdata (iCache_1_sram_1_ports_cmd_payload_wdata[511:0]  ), //i
    .sram_1_ports_cmd_payload_wstrb (iCache_1_sram_1_ports_cmd_payload_wstrb[63:0]   ), //i
    .sram_1_ports_rsp_valid         (sramBanks_2_sram_1_ports_rsp_valid              ), //o
    .sram_1_ports_rsp_payload_data  (sramBanks_2_sram_1_ports_rsp_payload_data[511:0]), //o
    .sram_2_ports_cmd_valid         (iCache_1_sram_2_ports_cmd_valid                 ), //i
    .sram_2_ports_cmd_payload_addr  (iCache_1_sram_2_ports_cmd_payload_addr[6:0]     ), //i
    .sram_2_ports_cmd_payload_wen   (iCache_1_sram_2_ports_cmd_payload_wen[15:0]     ), //i
    .sram_2_ports_cmd_payload_wdata (iCache_1_sram_2_ports_cmd_payload_wdata[511:0]  ), //i
    .sram_2_ports_cmd_payload_wstrb (iCache_1_sram_2_ports_cmd_payload_wstrb[63:0]   ), //i
    .sram_2_ports_rsp_valid         (sramBanks_2_sram_2_ports_rsp_valid              ), //o
    .sram_2_ports_rsp_payload_data  (sramBanks_2_sram_2_ports_rsp_payload_data[511:0]), //o
    .sram_3_ports_cmd_valid         (iCache_1_sram_3_ports_cmd_valid                 ), //i
    .sram_3_ports_cmd_payload_addr  (iCache_1_sram_3_ports_cmd_payload_addr[6:0]     ), //i
    .sram_3_ports_cmd_payload_wen   (iCache_1_sram_3_ports_cmd_payload_wen[15:0]     ), //i
    .sram_3_ports_cmd_payload_wdata (iCache_1_sram_3_ports_cmd_payload_wdata[511:0]  ), //i
    .sram_3_ports_cmd_payload_wstrb (iCache_1_sram_3_ports_cmd_payload_wstrb[63:0]   ), //i
    .sram_3_ports_rsp_valid         (sramBanks_2_sram_3_ports_rsp_valid              ), //o
    .sram_3_ports_rsp_payload_data  (sramBanks_2_sram_3_ports_rsp_payload_data[511:0]), //o
    .clk                            (clk                                             ), //i
    .reset                          (reset                                           )  //i
  );
  DCache dCache_1 (
    .stall                          (dCache_1_stall                                    ), //o
    .flush                          (1'b0                                              ), //i
    .cpu_cmd_valid                  (DCachePlugin_dcache_access_cmd_valid              ), //i
    .cpu_cmd_ready                  (dCache_1_cpu_cmd_ready                            ), //o
    .cpu_cmd_payload_addr           (DCachePlugin_dcache_access_cmd_payload_addr[63:0] ), //i
    .cpu_cmd_payload_wen            (DCachePlugin_dcache_access_cmd_payload_wen        ), //i
    .cpu_cmd_payload_wdata          (DCachePlugin_dcache_access_cmd_payload_wdata[63:0]), //i
    .cpu_cmd_payload_wstrb          (DCachePlugin_dcache_access_cmd_payload_wstrb[7:0] ), //i
    .cpu_rsp_valid                  (dCache_1_cpu_rsp_valid                            ), //o
    .cpu_rsp_payload_data           (dCache_1_cpu_rsp_payload_data[63:0]               ), //o
    .sram_0_ports_cmd_valid         (dCache_1_sram_0_ports_cmd_valid                   ), //o
    .sram_0_ports_cmd_payload_addr  (dCache_1_sram_0_ports_cmd_payload_addr[6:0]       ), //o
    .sram_0_ports_cmd_payload_wen   (dCache_1_sram_0_ports_cmd_payload_wen[7:0]        ), //o
    .sram_0_ports_cmd_payload_wdata (dCache_1_sram_0_ports_cmd_payload_wdata[511:0]    ), //o
    .sram_0_ports_cmd_payload_wstrb (dCache_1_sram_0_ports_cmd_payload_wstrb[63:0]     ), //o
    .sram_0_ports_rsp_valid         (sramBanks_3_sram_0_ports_rsp_valid                ), //i
    .sram_0_ports_rsp_payload_data  (sramBanks_3_sram_0_ports_rsp_payload_data[511:0]  ), //i
    .sram_1_ports_cmd_valid         (dCache_1_sram_1_ports_cmd_valid                   ), //o
    .sram_1_ports_cmd_payload_addr  (dCache_1_sram_1_ports_cmd_payload_addr[6:0]       ), //o
    .sram_1_ports_cmd_payload_wen   (dCache_1_sram_1_ports_cmd_payload_wen[7:0]        ), //o
    .sram_1_ports_cmd_payload_wdata (dCache_1_sram_1_ports_cmd_payload_wdata[511:0]    ), //o
    .sram_1_ports_cmd_payload_wstrb (dCache_1_sram_1_ports_cmd_payload_wstrb[63:0]     ), //o
    .sram_1_ports_rsp_valid         (sramBanks_3_sram_1_ports_rsp_valid                ), //i
    .sram_1_ports_rsp_payload_data  (sramBanks_3_sram_1_ports_rsp_payload_data[511:0]  ), //i
    .sram_2_ports_cmd_valid         (dCache_1_sram_2_ports_cmd_valid                   ), //o
    .sram_2_ports_cmd_payload_addr  (dCache_1_sram_2_ports_cmd_payload_addr[6:0]       ), //o
    .sram_2_ports_cmd_payload_wen   (dCache_1_sram_2_ports_cmd_payload_wen[7:0]        ), //o
    .sram_2_ports_cmd_payload_wdata (dCache_1_sram_2_ports_cmd_payload_wdata[511:0]    ), //o
    .sram_2_ports_cmd_payload_wstrb (dCache_1_sram_2_ports_cmd_payload_wstrb[63:0]     ), //o
    .sram_2_ports_rsp_valid         (sramBanks_3_sram_2_ports_rsp_valid                ), //i
    .sram_2_ports_rsp_payload_data  (sramBanks_3_sram_2_ports_rsp_payload_data[511:0]  ), //i
    .sram_3_ports_cmd_valid         (dCache_1_sram_3_ports_cmd_valid                   ), //o
    .sram_3_ports_cmd_payload_addr  (dCache_1_sram_3_ports_cmd_payload_addr[6:0]       ), //o
    .sram_3_ports_cmd_payload_wen   (dCache_1_sram_3_ports_cmd_payload_wen[7:0]        ), //o
    .sram_3_ports_cmd_payload_wdata (dCache_1_sram_3_ports_cmd_payload_wdata[511:0]    ), //o
    .sram_3_ports_cmd_payload_wstrb (dCache_1_sram_3_ports_cmd_payload_wstrb[63:0]     ), //o
    .sram_3_ports_rsp_valid         (sramBanks_3_sram_3_ports_rsp_valid                ), //i
    .sram_3_ports_rsp_payload_data  (sramBanks_3_sram_3_ports_rsp_payload_data[511:0]  ), //i
    .next_level_cmd_valid           (dCache_1_next_level_cmd_valid                     ), //o
    .next_level_cmd_ready           (dCache_1_next_level_cmd_ready                     ), //i
    .next_level_cmd_payload_addr    (dCache_1_next_level_cmd_payload_addr[63:0]        ), //o
    .next_level_cmd_payload_len     (dCache_1_next_level_cmd_payload_len[3:0]          ), //o
    .next_level_cmd_payload_size    (dCache_1_next_level_cmd_payload_size[2:0]         ), //o
    .next_level_cmd_payload_wen     (dCache_1_next_level_cmd_payload_wen               ), //o
    .next_level_cmd_payload_wdata   (dCache_1_next_level_cmd_payload_wdata[63:0]       ), //o
    .next_level_cmd_payload_wstrb   (dCache_1_next_level_cmd_payload_wstrb[7:0]        ), //o
    .next_level_rsp_valid           (dCache_1_next_level_rsp_valid                     ), //i
    .next_level_rsp_payload_data    (dcache_r_payload_data[63:0]                       ), //i
    .next_level_rsp_payload_bresp   (dcache_b_payload_resp[1:0]                        ), //i
    .next_level_rsp_payload_rvalid  (dcache_r_valid                                    ), //i
    .clk                            (clk                                               ), //i
    .reset                          (reset                                             )  //i
  );
  SramBanks_1 sramBanks_3 (
    .sram_0_ports_cmd_valid         (dCache_1_sram_0_ports_cmd_valid                 ), //i
    .sram_0_ports_cmd_payload_addr  (dCache_1_sram_0_ports_cmd_payload_addr[6:0]     ), //i
    .sram_0_ports_cmd_payload_wen   (dCache_1_sram_0_ports_cmd_payload_wen[7:0]      ), //i
    .sram_0_ports_cmd_payload_wdata (dCache_1_sram_0_ports_cmd_payload_wdata[511:0]  ), //i
    .sram_0_ports_cmd_payload_wstrb (dCache_1_sram_0_ports_cmd_payload_wstrb[63:0]   ), //i
    .sram_0_ports_rsp_valid         (sramBanks_3_sram_0_ports_rsp_valid              ), //o
    .sram_0_ports_rsp_payload_data  (sramBanks_3_sram_0_ports_rsp_payload_data[511:0]), //o
    .sram_1_ports_cmd_valid         (dCache_1_sram_1_ports_cmd_valid                 ), //i
    .sram_1_ports_cmd_payload_addr  (dCache_1_sram_1_ports_cmd_payload_addr[6:0]     ), //i
    .sram_1_ports_cmd_payload_wen   (dCache_1_sram_1_ports_cmd_payload_wen[7:0]      ), //i
    .sram_1_ports_cmd_payload_wdata (dCache_1_sram_1_ports_cmd_payload_wdata[511:0]  ), //i
    .sram_1_ports_cmd_payload_wstrb (dCache_1_sram_1_ports_cmd_payload_wstrb[63:0]   ), //i
    .sram_1_ports_rsp_valid         (sramBanks_3_sram_1_ports_rsp_valid              ), //o
    .sram_1_ports_rsp_payload_data  (sramBanks_3_sram_1_ports_rsp_payload_data[511:0]), //o
    .sram_2_ports_cmd_valid         (dCache_1_sram_2_ports_cmd_valid                 ), //i
    .sram_2_ports_cmd_payload_addr  (dCache_1_sram_2_ports_cmd_payload_addr[6:0]     ), //i
    .sram_2_ports_cmd_payload_wen   (dCache_1_sram_2_ports_cmd_payload_wen[7:0]      ), //i
    .sram_2_ports_cmd_payload_wdata (dCache_1_sram_2_ports_cmd_payload_wdata[511:0]  ), //i
    .sram_2_ports_cmd_payload_wstrb (dCache_1_sram_2_ports_cmd_payload_wstrb[63:0]   ), //i
    .sram_2_ports_rsp_valid         (sramBanks_3_sram_2_ports_rsp_valid              ), //o
    .sram_2_ports_rsp_payload_data  (sramBanks_3_sram_2_ports_rsp_payload_data[511:0]), //o
    .sram_3_ports_cmd_valid         (dCache_1_sram_3_ports_cmd_valid                 ), //i
    .sram_3_ports_cmd_payload_addr  (dCache_1_sram_3_ports_cmd_payload_addr[6:0]     ), //i
    .sram_3_ports_cmd_payload_wen   (dCache_1_sram_3_ports_cmd_payload_wen[7:0]      ), //i
    .sram_3_ports_cmd_payload_wdata (dCache_1_sram_3_ports_cmd_payload_wdata[511:0]  ), //i
    .sram_3_ports_cmd_payload_wstrb (dCache_1_sram_3_ports_cmd_payload_wstrb[63:0]   ), //i
    .sram_3_ports_rsp_valid         (sramBanks_3_sram_3_ports_rsp_valid              ), //o
    .sram_3_ports_rsp_payload_data  (sramBanks_3_sram_3_ports_rsp_payload_data[511:0]), //o
    .clk                            (clk                                             ), //i
    .reset                          (reset                                           )  //i
  );
  assign writeback_RD = (writeback_IS_LOAD ? writeback_LSU_RDATA : writeback_ALU_RESULT);
  assign memaccess_LSU_HOLD = DCachePlugin_dcache_access_stall;
  assign memaccess_TIMER_CEN = ((memaccess_LSUPlugin_is_timer && memaccess_LSUPlugin_is_mem) && memaccess_arbitration_isFiring);
  assign memaccess_LSU_WDATA = memaccess_LSUPlugin_lsu_wdata;
  assign execute_INT_HOLD = clint_1_int_hold;
  assign execute_REDIRECT_PC_NEXT = execute_ALUPlugin_redirect_pc_next;
  assign execute_REDIRECT_VALID = execute_ALUPlugin_redirect_valid;
  assign execute_IS_RET = execute_ALUPlugin_is_ret;
  assign execute_IS_CALL = execute_ALUPlugin_is_call;
  assign execute_IS_JMP = execute_ALUPlugin_is_jmp;
  assign execute_BRANCH_HISTORY = execute_ALUPlugin_branch_history;
  assign execute_BRANCH_TAKEN = execute_ALUPlugin_branch_taken;
  assign execute_BRANCH_OR_JUMP = (execute_ALUPlugin_branch_or_jump && execute_arbitration_isFiring);
  assign execute_BRANCH_OR_JALR = execute_ALUPlugin_branch_or_jalr;
  assign execute_MEM_WDATA = (execute_RS2_FROM_WB ? _zz_execute_MEM_WDATA_2 : (execute_RS2_FROM_MEM ? _zz_execute_MEM_WDATA_1 : (execute_RS2_FROM_LOAD ? _zz_execute_MEM_WDATA : execute_RS2)));
  assign execute_ALU_RESULT = execute_ALUPlugin_alu_result;
  assign decode_CSR_RDATA = csrRegfile_1_cpu_ports_rdata;
  assign execute_CSR_WEN = decode_to_execute_CSR_WEN;
  assign decode_CSR_WEN = decode_DecodePlugin_csr_wen;
  assign execute_CSR_ADDR = decode_to_execute_CSR_ADDR;
  assign decode_CSR_ADDR = decode_DecodePlugin_csr_addr;
  assign decode_CSR_CTRL = decode_DecodePlugin_csr_ctrl;
  assign execute_IS_STORE = decode_to_execute_IS_STORE;
  assign decode_IS_STORE = decode_DecodePlugin_is_store;
  assign execute_IS_LOAD = decode_to_execute_IS_LOAD;
  assign decode_IS_LOAD = decode_DecodePlugin_is_load;
  assign writeback_RD_ADDR = memaccess_to_writeback_RD_ADDR;
  assign memaccess_RD_ADDR = execute_to_memaccess_RD_ADDR;
  assign decode_RD_ADDR = decode_DecodePlugin_rd_addr;
  assign writeback_RD_WEN = memaccess_to_writeback_RD_WEN;
  assign memaccess_RD_WEN = execute_to_memaccess_RD_WEN;
  assign execute_RD_WEN = decode_to_execute_RD_WEN;
  assign decode_RD_WEN = decode_DecodePlugin_rd_wen;
  assign execute_MEM_CTRL = decode_to_execute_MEM_CTRL;
  assign decode_MEM_CTRL = decode_DecodePlugin_mem_ctrl;
  assign decode_SRC2_IS_IMM = decode_DecodePlugin_src2_is_imm;
  assign decode_ALU_WORD = decode_DecodePlugin_alu_word;
  assign decode_ALU_CTRL = decode_DecodePlugin_alu_ctrl;
  assign execute_RS2_ADDR = decode_to_execute_RS2_ADDR;
  assign decode_RS2_ADDR = decode_DecodePlugin_rs2_addr;
  assign decode_RS1_ADDR = decode_DecodePlugin_rs1_addr;
  assign decode_RS2 = decode_DecodePlugin_rs2;
  assign decode_RS1 = decode_DecodePlugin_rs1;
  assign decode_IMM = decode_DecodePlugin_imm;
  assign fetch_INT_PC = clint_1_int_pc;
  assign fetch_INT_EN = clint_1_int_en;
  assign fetch_PREDICT_PC = pc_next;
  assign decode_PREDICT_TAKEN = fetch_to_decode_PREDICT_TAKEN;
  assign fetch_PREDICT_TAKEN = fetch_FetchPlugin_predict_taken_out_payload;
  assign fetch_PREDICT_VALID = ICachePlugin_icache_access_cmd_fire_4;
  assign memaccess_INSTRUCTION = execute_to_memaccess_INSTRUCTION;
  assign execute_INSTRUCTION = decode_to_execute_INSTRUCTION;
  assign fetch_INSTRUCTION = fetch_FetchPlugin_instruction_out_stream_payload;
  assign decode_PC_NEXT = fetch_to_decode_PC_NEXT;
  assign fetch_PC_NEXT = fetch_FetchPlugin_pc_stream_fifo_next_payload;
  assign memaccess_PC = execute_to_memaccess_PC;
  assign fetch_PC = fetch_FetchPlugin_pc_out_stream_payload;
  assign writeback_INSTRUCTION = memaccess_to_writeback_INSTRUCTION;
  assign writeback_PC = memaccess_to_writeback_PC;
  assign writeback_ALU_RESULT = memaccess_to_writeback_ALU_RESULT;
  assign writeback_LSU_RDATA = memaccess_to_writeback_LSU_RDATA;
  assign writeback_IS_LOAD = memaccess_to_writeback_IS_LOAD;
  assign memaccess_MEM_CTRL = execute_to_memaccess_MEM_CTRL;
  assign memaccess_MEM_WDATA = execute_to_memaccess_MEM_WDATA;
  assign memaccess_IS_STORE = execute_to_memaccess_IS_STORE;
  assign memaccess_IS_LOAD = execute_to_memaccess_IS_LOAD;
  assign execute_CSR_CTRL = decode_to_execute_CSR_CTRL;
  assign execute_SRC1 = execute_ALUPlugin_src1;
  assign _zz_ecall = execute_CSR_CTRL;
  assign _zz_decode_to_execute_CSR_ADDR = decode_CSR_ADDR;
  assign _zz_memaccess_arbitration_haltItself = memaccess_LSU_HOLD;
  assign _zz_DecodePlugin_hazard_ctrl_rs1_from_mem = execute_BRANCH_OR_JALR;
  assign _zz_DecodePlugin_hazard_rs2_from_mem = execute_RS2_ADDR;
  assign _zz_DecodePlugin_hazard_rs1_from_mem = memaccess_IS_LOAD;
  assign _zz_DecodePlugin_hazard_rs1_from_mem_1 = execute_RS1_ADDR;
  assign _zz_DecodePlugin_hazard_rs1_from_mem_2 = memaccess_RD_ADDR;
  assign _zz_DecodePlugin_hazard_rs1_from_mem_3 = memaccess_RD_WEN;
  assign execute_PC_NEXT = decode_to_execute_PC_NEXT;
  assign execute_PREDICT_TAKEN = decode_to_execute_PREDICT_TAKEN;
  assign execute_CSR_RDATA = decode_to_execute_CSR_RDATA;
  assign execute_ALU_WORD = decode_to_execute_ALU_WORD;
  assign execute_CTRL_RS2_FROM_WB = DecodePlugin_hazard_ctrl_rs2_from_wb;
  assign execute_CTRL_RS2_FROM_LOAD = DecodePlugin_hazard_ctrl_rs2_from_load;
  assign execute_CTRL_RS2_FROM_MEM = DecodePlugin_hazard_ctrl_rs2_from_mem;
  assign execute_CTRL_RS1_FROM_WB = DecodePlugin_hazard_ctrl_rs1_from_wb;
  assign _zz_execute_MEM_WDATA = memaccess_LSU_RDATA;
  assign execute_CTRL_RS1_FROM_LOAD = DecodePlugin_hazard_ctrl_rs1_from_load;
  assign _zz_execute_MEM_WDATA_1 = memaccess_ALU_RESULT;
  assign execute_CTRL_RS1_FROM_MEM = DecodePlugin_hazard_ctrl_rs1_from_mem;
  assign execute_RS2 = decode_to_execute_RS2;
  assign execute_RS2_FROM_WB = DecodePlugin_hazard_rs2_from_wb;
  assign execute_RS2_FROM_LOAD = DecodePlugin_hazard_rs2_from_load;
  assign execute_RS2_FROM_MEM = DecodePlugin_hazard_rs2_from_mem;
  assign execute_IMM = decode_to_execute_IMM;
  assign execute_SRC2_IS_IMM = decode_to_execute_SRC2_IS_IMM;
  assign execute_RS1 = decode_to_execute_RS1;
  assign execute_RS1_FROM_WB = DecodePlugin_hazard_rs1_from_wb;
  assign memaccess_LSU_RDATA = memaccess_LSUPlugin_lsu_rdata;
  assign execute_RS1_FROM_LOAD = DecodePlugin_hazard_rs1_from_load;
  assign memaccess_ALU_RESULT = execute_to_memaccess_ALU_RESULT;
  assign execute_RS1_FROM_MEM = DecodePlugin_hazard_rs1_from_mem;
  assign execute_PC = decode_to_execute_PC;
  assign execute_RS1_ADDR = decode_to_execute_RS1_ADDR;
  assign execute_RD_ADDR = decode_to_execute_RD_ADDR;
  assign execute_ALU_CTRL = decode_to_execute_ALU_CTRL;
  assign _zz_execute_MEM_WDATA_2 = writeback_RD;
  assign _zz_DecodePlugin_hazard_rs1_from_wb = writeback_RD_ADDR;
  assign _zz_DecodePlugin_hazard_rs1_from_wb_1 = writeback_RD_WEN;
  assign decode_INSTRUCTION = fetch_to_decode_INSTRUCTION;
  assign decode_PC = fetch_to_decode_PC;
  assign _zz_execute_to_memaccess_PC = execute_PC;
  assign fetch_BPU_PC_NEXT = gshare_predictor_1_predict_pc_next;
  assign _zz_pc_next = execute_REDIRECT_PC_NEXT;
  assign when_FetchPlugin_l97 = execute_REDIRECT_VALID;
  assign fetch_BPU_BRANCH_TAKEN = gshare_predictor_1_predict_taken;
  assign when_FetchPlugin_l94 = fetch_INT_EN;
  assign fetch_arbitration_haltByOther = 1'b0;
  always @(*) begin
    fetch_arbitration_removeIt = 1'b0;
    if(fetch_arbitration_isFlushed) begin
      fetch_arbitration_removeIt = 1'b1;
    end
  end

  assign fetch_arbitration_flushNext = 1'b0;
  assign decode_arbitration_haltByOther = 1'b0;
  always @(*) begin
    decode_arbitration_removeIt = 1'b0;
    if(decode_arbitration_isFlushed) begin
      decode_arbitration_removeIt = 1'b1;
    end
  end

  assign decode_arbitration_flushNext = 1'b0;
  assign execute_arbitration_haltByOther = 1'b0;
  always @(*) begin
    execute_arbitration_removeIt = 1'b0;
    if(execute_arbitration_isFlushed) begin
      execute_arbitration_removeIt = 1'b1;
    end
  end

  assign execute_arbitration_flushNext = 1'b0;
  assign memaccess_arbitration_haltByOther = 1'b0;
  always @(*) begin
    memaccess_arbitration_removeIt = 1'b0;
    if(memaccess_arbitration_isFlushed) begin
      memaccess_arbitration_removeIt = 1'b1;
    end
  end

  assign memaccess_arbitration_flushNext = 1'b0;
  assign writeback_arbitration_haltByOther = 1'b0;
  always @(*) begin
    writeback_arbitration_removeIt = 1'b0;
    if(writeback_arbitration_isFlushed) begin
      writeback_arbitration_removeIt = 1'b1;
    end
  end

  assign writeback_arbitration_flushNext = 1'b0;
  assign fetch_FetchPlugin_fetch_flush = (when_FetchPlugin_l94 || fetch_arbitration_flushIt);
  assign ICachePlugin_icache_access_cmd_fire = (ICachePlugin_icache_access_cmd_valid && ICachePlugin_icache_access_cmd_ready);
  assign fetch_FetchPlugin_bpu_predict_taken = (fetch_BPU_BRANCH_TAKEN && ICachePlugin_icache_access_cmd_fire);
  assign fetch_FetchPlugin_fifo_all_valid = ((fetch_FetchPlugin_pc_out_stream_valid && fetch_FetchPlugin_instruction_out_stream_valid) && fetch_FetchPlugin_pc_stream_fifo_next_valid);
  assign IDLE = 2'b00;
  assign FETCH = 2'b01;
  assign HALT = 2'b11;
  assign when_FetchPlugin_l64 = (! fetch_arbitration_isStuck);
  always @(*) begin
    if((fetch_state == IDLE)) begin
        if(when_FetchPlugin_l64) begin
          fetch_state_next = FETCH;
        end else begin
          fetch_state_next = IDLE;
        end
    end else if((fetch_state == FETCH)) begin
        if(when_FetchPlugin_l72) begin
          fetch_state_next = HALT;
        end else begin
          fetch_state_next = FETCH;
        end
    end else if((fetch_state == HALT)) begin
        if(when_FetchPlugin_l80) begin
          fetch_state_next = FETCH;
        end else begin
          fetch_state_next = HALT;
        end
    end else begin
        fetch_state_next = IDLE;
    end
  end

  assign ICachePlugin_icache_access_cmd_isStall = (ICachePlugin_icache_access_cmd_valid && (! ICachePlugin_icache_access_cmd_ready));
  assign when_FetchPlugin_l72 = (ICachePlugin_icache_access_cmd_isStall || fetch_arbitration_isStuck);
  assign when_FetchPlugin_l80 = (ICachePlugin_icache_access_cmd_ready && (! fetch_arbitration_isStuck));
  assign when_FetchPlugin_l93 = (! ICachePlugin_icache_access_cmd_ready);
  assign when_FetchPlugin_l109 = (fetch_state_next == FETCH);
  assign ICachePlugin_icache_access_cmd_fire_1 = (ICachePlugin_icache_access_cmd_valid && ICachePlugin_icache_access_cmd_ready);
  assign ICachePlugin_icache_access_cmd_fire_2 = (ICachePlugin_icache_access_cmd_valid && ICachePlugin_icache_access_cmd_ready);
  assign fetch_FetchPlugin_pc_in_stream_valid = ICachePlugin_icache_access_cmd_fire_2;
  assign fetch_FetchPlugin_pc_in_stream_payload = pc_next;
  assign fetch_FetchPlugin_pc_out_stream_ready = fetch_arbitration_isFiring;
  assign fetch_FetchPlugin_pc_in_stream_ready = fetch_FetchPlugin_pc_stream_fifo_ports_s_ports_ready;
  assign fetch_FetchPlugin_pc_out_stream_valid = fetch_FetchPlugin_pc_stream_fifo_ports_m_ports_valid;
  assign fetch_FetchPlugin_pc_out_stream_payload = fetch_FetchPlugin_pc_stream_fifo_ports_m_ports_payload;
  assign ICachePlugin_icache_access_cmd_fire_3 = (ICachePlugin_icache_access_cmd_valid && ICachePlugin_icache_access_cmd_ready);
  assign fetch_FetchPlugin_predict_taken_in_valid = ICachePlugin_icache_access_cmd_fire_3;
  assign fetch_FetchPlugin_predict_taken_in_payload = fetch_BPU_BRANCH_TAKEN;
  assign fetch_FetchPlugin_predict_taken_out_ready = fetch_arbitration_isFiring;
  assign fetch_FetchPlugin_predict_taken_in_ready = fetch_FetchPlugin_predict_taken_fifo_ports_s_ports_ready;
  assign fetch_FetchPlugin_predict_taken_out_valid = fetch_FetchPlugin_predict_taken_fifo_ports_m_ports_valid;
  assign fetch_FetchPlugin_predict_taken_out_payload = fetch_FetchPlugin_predict_taken_fifo_ports_m_ports_payload;
  assign fetch_FetchPlugin_instruction_in_stream_valid = ((ICachePlugin_icache_access_rsp_valid && (! rsp_flush)) && (! fetch_FetchPlugin_fetch_flush));
  assign fetch_FetchPlugin_instruction_in_stream_payload = ICachePlugin_icache_access_rsp_payload_data;
  assign fetch_FetchPlugin_instruction_out_stream_ready = fetch_arbitration_isFiring;
  assign fetch_FetchPlugin_instruction_in_stream_ready = fetch_FetchPlugin_instruction_stream_fifo_ports_s_ports_ready;
  assign fetch_FetchPlugin_instruction_out_stream_valid = fetch_FetchPlugin_instruction_stream_fifo_ports_m_ports_valid;
  assign fetch_FetchPlugin_instruction_out_stream_payload = fetch_FetchPlugin_instruction_stream_fifo_ports_m_ports_payload;
  assign ICachePlugin_icache_access_cmd_fire_4 = (ICachePlugin_icache_access_cmd_valid && ICachePlugin_icache_access_cmd_ready);
  assign fetch_arbitration_isValid = ((fetch_FetchPlugin_fifo_all_valid && (! fetch_arbitration_isStuck)) && (! fetch_FetchPlugin_fetch_flush));
  assign ICachePlugin_icache_access_cmd_valid = (fetch_valid && (! fetch_FetchPlugin_fetch_flush));
  assign ICachePlugin_icache_access_cmd_payload_addr = pc_next;
  assign decode_DecodePlugin_rs1_req = (! (((decode_INSTRUCTION[6 : 0] == 7'h37) || (decode_INSTRUCTION[6 : 0] == 7'h17)) || (decode_INSTRUCTION[6 : 0] == 7'h6f)));
  assign decode_DecodePlugin_rs2_req = (! ((((decode_INSTRUCTION[6 : 0] == 7'h37) || (decode_INSTRUCTION[6 : 0] == 7'h17)) || (decode_INSTRUCTION[6 : 0] == 7'h6f)) || ((((decode_INSTRUCTION[6 : 0] == 7'h13) || (decode_INSTRUCTION[6 : 0] == 7'h1b)) || (decode_INSTRUCTION[6 : 0] == 7'h03)) || (decode_INSTRUCTION[6 : 0] == 7'h67))));
  assign decode_DecodePlugin_rs1_addr = decode_INSTRUCTION[19 : 15];
  assign decode_DecodePlugin_rs2_addr = decode_INSTRUCTION[24 : 20];
  assign decode_DecodePlugin_rd_addr = decode_INSTRUCTION[11 : 7];
  assign decode_DecodePlugin_alu_word = ((decode_INSTRUCTION[6 : 0] == 7'h3b) || (decode_INSTRUCTION[6 : 0] == 7'h1b));
  assign decode_DecodePlugin_src2_is_imm = ((((((decode_INSTRUCTION[6 : 0] == 7'h13) || (decode_INSTRUCTION[6 : 0] == 7'h1b)) || (decode_INSTRUCTION[6 : 0] == 7'h03)) || (decode_INSTRUCTION[6 : 0] == 7'h67)) || (decode_INSTRUCTION[6 : 0] == 7'h23)) || ((decode_INSTRUCTION[6 : 0] == 7'h37) || (decode_INSTRUCTION[6 : 0] == 7'h17)));
  assign decode_DecodePlugin_csr_addr = decode_INSTRUCTION[31 : 20];
  assign decode_DecodePlugin_csr_wen = (((decode_DecodePlugin_csr_ctrl == CsrCtrlEnum_CSRRW) || (decode_DecodePlugin_csr_ctrl == CsrCtrlEnum_CSRRS)) || (decode_DecodePlugin_csr_ctrl == CsrCtrlEnum_CSRRC));
  assign when_DecodePlugin_l116 = ((((decode_INSTRUCTION[6 : 0] == 7'h13) || (decode_INSTRUCTION[6 : 0] == 7'h1b)) || (decode_INSTRUCTION[6 : 0] == 7'h03)) || (decode_INSTRUCTION[6 : 0] == 7'h67));
  assign _zz_decode_DecodePlugin_imm = decode_INSTRUCTION[31];
  always @(*) begin
    _zz_decode_DecodePlugin_imm_1[51] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[50] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[49] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[48] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[47] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[46] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[45] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[44] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[43] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[42] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[41] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[40] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[39] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[38] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[37] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[36] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[35] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[34] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[33] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[32] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[31] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[30] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[29] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[28] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[27] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[26] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[25] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[24] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[23] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[22] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[21] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[20] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[19] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[18] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[17] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[16] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[15] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[14] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[13] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[12] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[11] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[10] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[9] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[8] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[7] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[6] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[5] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[4] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[3] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[2] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[1] = _zz_decode_DecodePlugin_imm;
    _zz_decode_DecodePlugin_imm_1[0] = _zz_decode_DecodePlugin_imm;
  end

  always @(*) begin
    if(when_DecodePlugin_l116) begin
      decode_DecodePlugin_imm = {_zz_decode_DecodePlugin_imm_1,decode_INSTRUCTION[31 : 20]};
    end else begin
      if(when_DecodePlugin_l119) begin
        decode_DecodePlugin_imm = {_zz_decode_DecodePlugin_imm_3,{decode_INSTRUCTION[31 : 25],decode_INSTRUCTION[11 : 7]}};
      end else begin
        if(when_DecodePlugin_l122) begin
          decode_DecodePlugin_imm = {{_zz_decode_DecodePlugin_imm_5,{{{decode_INSTRUCTION[31],decode_INSTRUCTION[7]},decode_INSTRUCTION[30 : 25]},decode_INSTRUCTION[11 : 8]}},1'b0};
        end else begin
          if(when_DecodePlugin_l125) begin
            decode_DecodePlugin_imm = {{_zz_decode_DecodePlugin_imm_7,{{{decode_INSTRUCTION[31],decode_INSTRUCTION[19 : 12]},decode_INSTRUCTION[20]},decode_INSTRUCTION[30 : 21]}},1'b0};
          end else begin
            if(when_DecodePlugin_l128) begin
              decode_DecodePlugin_imm = {_zz_decode_DecodePlugin_imm_9,{decode_INSTRUCTION[31 : 12],12'h0}};
            end else begin
              decode_DecodePlugin_imm = {_zz_decode_DecodePlugin_imm_11,decode_INSTRUCTION[31 : 20]};
            end
          end
        end
      end
    end
  end

  assign _zz_decode_DecodePlugin_imm_2 = _zz__zz_decode_DecodePlugin_imm_2[11];
  always @(*) begin
    _zz_decode_DecodePlugin_imm_3[51] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[50] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[49] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[48] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[47] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[46] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[45] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[44] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[43] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[42] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[41] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[40] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[39] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[38] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[37] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[36] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[35] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[34] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[33] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[32] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[31] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[30] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[29] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[28] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[27] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[26] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[25] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[24] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[23] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[22] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[21] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[20] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[19] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[18] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[17] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[16] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[15] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[14] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[13] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[12] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[11] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[10] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[9] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[8] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[7] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[6] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[5] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[4] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[3] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[2] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[1] = _zz_decode_DecodePlugin_imm_2;
    _zz_decode_DecodePlugin_imm_3[0] = _zz_decode_DecodePlugin_imm_2;
  end

  assign _zz_decode_DecodePlugin_imm_4 = _zz__zz_decode_DecodePlugin_imm_4[11];
  always @(*) begin
    _zz_decode_DecodePlugin_imm_5[50] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[49] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[48] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[47] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[46] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[45] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[44] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[43] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[42] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[41] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[40] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[39] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[38] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[37] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[36] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[35] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[34] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[33] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[32] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[31] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[30] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[29] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[28] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[27] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[26] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[25] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[24] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[23] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[22] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[21] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[20] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[19] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[18] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[17] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[16] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[15] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[14] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[13] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[12] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[11] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[10] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[9] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[8] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[7] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[6] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[5] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[4] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[3] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[2] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[1] = _zz_decode_DecodePlugin_imm_4;
    _zz_decode_DecodePlugin_imm_5[0] = _zz_decode_DecodePlugin_imm_4;
  end

  assign _zz_decode_DecodePlugin_imm_6 = _zz__zz_decode_DecodePlugin_imm_6[19];
  always @(*) begin
    _zz_decode_DecodePlugin_imm_7[42] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[41] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[40] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[39] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[38] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[37] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[36] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[35] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[34] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[33] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[32] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[31] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[30] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[29] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[28] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[27] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[26] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[25] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[24] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[23] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[22] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[21] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[20] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[19] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[18] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[17] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[16] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[15] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[14] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[13] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[12] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[11] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[10] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[9] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[8] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[7] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[6] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[5] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[4] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[3] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[2] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[1] = _zz_decode_DecodePlugin_imm_6;
    _zz_decode_DecodePlugin_imm_7[0] = _zz_decode_DecodePlugin_imm_6;
  end

  assign _zz_decode_DecodePlugin_imm_8 = _zz__zz_decode_DecodePlugin_imm_8[31];
  always @(*) begin
    _zz_decode_DecodePlugin_imm_9[31] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[30] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[29] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[28] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[27] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[26] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[25] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[24] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[23] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[22] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[21] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[20] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[19] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[18] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[17] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[16] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[15] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[14] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[13] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[12] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[11] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[10] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[9] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[8] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[7] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[6] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[5] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[4] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[3] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[2] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[1] = _zz_decode_DecodePlugin_imm_8;
    _zz_decode_DecodePlugin_imm_9[0] = _zz_decode_DecodePlugin_imm_8;
  end

  assign _zz_decode_DecodePlugin_imm_10 = decode_INSTRUCTION[31];
  always @(*) begin
    _zz_decode_DecodePlugin_imm_11[51] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[50] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[49] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[48] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[47] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[46] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[45] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[44] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[43] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[42] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[41] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[40] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[39] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[38] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[37] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[36] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[35] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[34] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[33] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[32] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[31] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[30] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[29] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[28] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[27] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[26] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[25] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[24] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[23] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[22] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[21] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[20] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[19] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[18] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[17] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[16] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[15] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[14] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[13] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[12] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[11] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[10] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[9] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[8] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[7] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[6] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[5] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[4] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[3] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[2] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[1] = _zz_decode_DecodePlugin_imm_10;
    _zz_decode_DecodePlugin_imm_11[0] = _zz_decode_DecodePlugin_imm_10;
  end

  assign when_DecodePlugin_l119 = (decode_INSTRUCTION[6 : 0] == 7'h23);
  assign when_DecodePlugin_l122 = (decode_INSTRUCTION[6 : 0] == 7'h63);
  assign when_DecodePlugin_l125 = (decode_INSTRUCTION[6 : 0] == 7'h6f);
  assign when_DecodePlugin_l128 = ((decode_INSTRUCTION[6 : 0] == 7'h37) || (decode_INSTRUCTION[6 : 0] == 7'h17));
  always @(*) begin
    casez(decode_INSTRUCTION)
      32'b0000000??????????000?????0110011, 32'b0000000??????????000?????0111011, 32'b?????????????????000?????0010011, 32'b?????????????????000?????0011011, 32'b?????????????????000?????0100011, 32'b?????????????????001?????0100011, 32'b?????????????????010?????0100011, 32'b?????????????????011?????0100011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_ADD;
      end
      32'b0100000??????????000?????0110011, 32'b0100000??????????000?????0111011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_SUB;
      end
      32'b0000000??????????010?????0110011, 32'b?????????????????010?????0010011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_SLT;
      end
      32'b0000000??????????011?????0110011, 32'b?????????????????011?????0010011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_SLTU;
      end
      32'b0000000??????????100?????0110011, 32'b?????????????????100?????0010011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_XOR_1;
      end
      32'b0000000??????????001?????0110011, 32'b000000???????????001?????0010011, 32'b0000000??????????001?????0111011, 32'b000000???????????001?????0011011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_SLL_1;
      end
      32'b0000000??????????101?????0110011, 32'b000000???????????101?????0010011, 32'b0000000??????????101?????0111011, 32'b000000???????????101?????0011011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_SRL_1;
      end
      32'b0100000??????????101?????0110011, 32'b010000???????????101?????0010011, 32'b0100000??????????101?????0111011, 32'b010000???????????101?????0011011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_SRA_1;
      end
      32'b0000000??????????111?????0110011, 32'b?????????????????111?????0010011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_AND_1;
      end
      32'b0000000??????????110?????0110011, 32'b?????????????????110?????0010011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_OR_1;
      end
      32'b?????????????????????????0110111 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_LUI;
      end
      32'b?????????????????????????0010111 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_AUIPC;
      end
      32'b??????????0??????????????1101111 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_JAL;
      end
      32'b?????????????????000?????1100111 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_JALR;
      end
      32'b?????????????????000???0?1100011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_BEQ;
      end
      32'b?????????????????001???0?1100011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_BNE;
      end
      32'b?????????????????100???0?1100011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_BLT;
      end
      32'b?????????????????101???0?1100011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_BGE;
      end
      32'b?????????????????110???0?1100011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_BLTU;
      end
      32'b?????????????????111???0?1100011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_BGEU;
      end
      32'b?????????????????001?????1110011, 32'b?????????????????010?????1110011, 32'b?????????????????011?????1110011, 32'b?????????????????101?????1110011, 32'b?????????????????110?????1110011, 32'b?????????????????111?????1110011 : begin
        decode_DecodePlugin_alu_ctrl = AluCtrlEnum_CSR;
      end
      default : begin
        decode_DecodePlugin_alu_ctrl = 5'h0;
      end
    endcase
  end

  always @(*) begin
    casez(decode_INSTRUCTION)
      32'b?????????????????000?????0000011 : begin
        decode_DecodePlugin_mem_ctrl = MemCtrlEnum_LB;
      end
      32'b?????????????????100?????0000011 : begin
        decode_DecodePlugin_mem_ctrl = MemCtrlEnum_LBU;
      end
      32'b?????????????????001?????0000011 : begin
        decode_DecodePlugin_mem_ctrl = MemCtrlEnum_LH;
      end
      32'b?????????????????101?????0000011 : begin
        decode_DecodePlugin_mem_ctrl = MemCtrlEnum_LHU;
      end
      32'b?????????????????010?????0000011 : begin
        decode_DecodePlugin_mem_ctrl = MemCtrlEnum_LW;
      end
      32'b?????????????????110?????0000011 : begin
        decode_DecodePlugin_mem_ctrl = MemCtrlEnum_LWU;
      end
      32'b?????????????????011?????0000011 : begin
        decode_DecodePlugin_mem_ctrl = MemCtrlEnum_LD;
      end
      32'b?????????????????000?????0100011 : begin
        decode_DecodePlugin_mem_ctrl = MemCtrlEnum_SB;
      end
      32'b?????????????????001?????0100011 : begin
        decode_DecodePlugin_mem_ctrl = MemCtrlEnum_SH;
      end
      32'b?????????????????010?????0100011 : begin
        decode_DecodePlugin_mem_ctrl = MemCtrlEnum_SW;
      end
      32'b?????????????????011?????0100011 : begin
        decode_DecodePlugin_mem_ctrl = MemCtrlEnum_SD;
      end
      default : begin
        decode_DecodePlugin_mem_ctrl = 4'b0000;
      end
    endcase
  end

  always @(*) begin
    casez(decode_INSTRUCTION)
      32'b?????????????????000?????0000011 : begin
        decode_DecodePlugin_is_load = 1'b1;
      end
      32'b?????????????????100?????0000011 : begin
        decode_DecodePlugin_is_load = 1'b1;
      end
      32'b?????????????????001?????0000011 : begin
        decode_DecodePlugin_is_load = 1'b1;
      end
      32'b?????????????????101?????0000011 : begin
        decode_DecodePlugin_is_load = 1'b1;
      end
      32'b?????????????????010?????0000011 : begin
        decode_DecodePlugin_is_load = 1'b1;
      end
      32'b?????????????????110?????0000011 : begin
        decode_DecodePlugin_is_load = 1'b1;
      end
      32'b?????????????????011?????0000011 : begin
        decode_DecodePlugin_is_load = 1'b1;
      end
      32'b?????????????????000?????0100011 : begin
        decode_DecodePlugin_is_load = 1'b0;
      end
      32'b?????????????????001?????0100011 : begin
        decode_DecodePlugin_is_load = 1'b0;
      end
      32'b?????????????????010?????0100011 : begin
        decode_DecodePlugin_is_load = 1'b0;
      end
      32'b?????????????????011?????0100011 : begin
        decode_DecodePlugin_is_load = 1'b0;
      end
      default : begin
        decode_DecodePlugin_is_load = 1'b0;
      end
    endcase
  end

  always @(*) begin
    casez(decode_INSTRUCTION)
      32'b?????????????????000?????0000011 : begin
        decode_DecodePlugin_is_store = 1'b0;
      end
      32'b?????????????????100?????0000011 : begin
        decode_DecodePlugin_is_store = 1'b0;
      end
      32'b?????????????????001?????0000011 : begin
        decode_DecodePlugin_is_store = 1'b0;
      end
      32'b?????????????????101?????0000011 : begin
        decode_DecodePlugin_is_store = 1'b0;
      end
      32'b?????????????????010?????0000011 : begin
        decode_DecodePlugin_is_store = 1'b0;
      end
      32'b?????????????????110?????0000011 : begin
        decode_DecodePlugin_is_store = 1'b0;
      end
      32'b?????????????????011?????0000011 : begin
        decode_DecodePlugin_is_store = 1'b0;
      end
      32'b?????????????????000?????0100011 : begin
        decode_DecodePlugin_is_store = 1'b1;
      end
      32'b?????????????????001?????0100011 : begin
        decode_DecodePlugin_is_store = 1'b1;
      end
      32'b?????????????????010?????0100011 : begin
        decode_DecodePlugin_is_store = 1'b1;
      end
      32'b?????????????????011?????0100011 : begin
        decode_DecodePlugin_is_store = 1'b1;
      end
      default : begin
        decode_DecodePlugin_is_store = 1'b0;
      end
    endcase
  end

  always @(*) begin
    casez(decode_INSTRUCTION)
      32'b00000000000000000000000001110011 : begin
        decode_DecodePlugin_csr_ctrl = CsrCtrlEnum_ECALL;
      end
      32'b00000000000100000000000001110011 : begin
        decode_DecodePlugin_csr_ctrl = CsrCtrlEnum_EBREAK;
      end
      32'b00110000001000000000000001110011 : begin
        decode_DecodePlugin_csr_ctrl = CsrCtrlEnum_MRET;
      end
      32'b?????????????????001?????1110011 : begin
        decode_DecodePlugin_csr_ctrl = CsrCtrlEnum_CSRRW;
      end
      32'b?????????????????010?????1110011 : begin
        decode_DecodePlugin_csr_ctrl = CsrCtrlEnum_CSRRS;
      end
      32'b?????????????????011?????1110011 : begin
        decode_DecodePlugin_csr_ctrl = CsrCtrlEnum_CSRRC;
      end
      32'b?????????????????101?????1110011 : begin
        decode_DecodePlugin_csr_ctrl = CsrCtrlEnum_CSRRWI;
      end
      32'b?????????????????110?????1110011 : begin
        decode_DecodePlugin_csr_ctrl = CsrCtrlEnum_CSRRSI;
      end
      32'b?????????????????111?????1110011 : begin
        decode_DecodePlugin_csr_ctrl = CsrCtrlEnum_CSRRCI;
      end
      default : begin
        decode_DecodePlugin_csr_ctrl = 4'b0000;
      end
    endcase
  end

  assign decode_DecodePlugin_rs1 = regFileModule_1_read_ports_rs1_value;
  assign decode_DecodePlugin_rs2 = regFileModule_1_read_ports_rs2_value;
  assign decode_DecodePlugin_rd_wen = ((((((! (decode_INSTRUCTION[6 : 0] == 7'h23)) && (! (decode_INSTRUCTION[6 : 0] == 7'h63))) && (! ((decode_INSTRUCTION & 32'hffffffff) == 32'h00100073))) && (! ((decode_INSTRUCTION & 32'hffffffff) == 32'h00000073))) && (! ((decode_INSTRUCTION & 32'hffffffff) == 32'h30200073))) && (decode_INSTRUCTION[6 : 0] != 7'h0f));
  assign DecodePlugin_hazard_decode_rs1_req = decode_DecodePlugin_rs1_req;
  assign DecodePlugin_hazard_decode_rs2_req = decode_DecodePlugin_rs2_req;
  assign DecodePlugin_hazard_decode_rs1_addr = decode_DecodePlugin_rs1_addr;
  assign DecodePlugin_hazard_decode_rs2_addr = decode_DecodePlugin_rs2_addr;
  assign regFileModule_1_write_ports_rd_wen = (writeback_arbitration_isFiring && _zz_DecodePlugin_hazard_rs1_from_wb_1);
  assign execute_ALUPlugin_src1_word = execute_ALUPlugin_src1[31 : 0];
  assign execute_ALUPlugin_src2_word = execute_ALUPlugin_src2[31 : 0];
  assign execute_ALUPlugin_shift_bits = execute_ALUPlugin_src2[5 : 0];
  assign execute_ALUPlugin_add_result = ($signed(_zz_execute_ALUPlugin_add_result) + $signed(_zz_execute_ALUPlugin_add_result_1));
  assign execute_ALUPlugin_sub_result = ($signed(_zz_execute_ALUPlugin_sub_result) - $signed(_zz_execute_ALUPlugin_sub_result_1));
  assign execute_ALUPlugin_slt_result = ($signed(_zz_execute_ALUPlugin_slt_result) < $signed(_zz_execute_ALUPlugin_slt_result_1));
  assign execute_ALUPlugin_sltu_result = (execute_ALUPlugin_src1 < execute_ALUPlugin_src2);
  assign execute_ALUPlugin_xor_result = (execute_ALUPlugin_src1 ^ execute_ALUPlugin_src2);
  assign execute_ALUPlugin_sll_result = (execute_ALUPlugin_src1 <<< execute_ALUPlugin_shift_bits);
  assign execute_ALUPlugin_srl_result = (execute_ALUPlugin_src1 >>> execute_ALUPlugin_shift_bits);
  assign execute_ALUPlugin_sra_result = ($signed(_zz_execute_ALUPlugin_sra_result) >>> execute_ALUPlugin_shift_bits);
  assign execute_ALUPlugin_and_result = (execute_ALUPlugin_src1 & execute_ALUPlugin_src2);
  assign execute_ALUPlugin_or_result = (execute_ALUPlugin_src1 | execute_ALUPlugin_src2);
  assign _zz_execute_ALUPlugin_addw_result = execute_ALUPlugin_add_result[31];
  always @(*) begin
    _zz_execute_ALUPlugin_addw_result_1[31] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[30] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[29] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[28] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[27] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[26] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[25] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[24] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[23] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[22] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[21] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[20] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[19] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[18] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[17] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[16] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[15] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[14] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[13] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[12] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[11] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[10] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[9] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[8] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[7] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[6] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[5] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[4] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[3] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[2] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[1] = _zz_execute_ALUPlugin_addw_result;
    _zz_execute_ALUPlugin_addw_result_1[0] = _zz_execute_ALUPlugin_addw_result;
  end

  assign execute_ALUPlugin_addw_result = {_zz_execute_ALUPlugin_addw_result_1,_zz_execute_ALUPlugin_addw_result_2};
  assign _zz_execute_ALUPlugin_subw_result = execute_ALUPlugin_sub_result[31];
  always @(*) begin
    _zz_execute_ALUPlugin_subw_result_1[31] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[30] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[29] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[28] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[27] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[26] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[25] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[24] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[23] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[22] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[21] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[20] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[19] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[18] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[17] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[16] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[15] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[14] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[13] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[12] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[11] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[10] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[9] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[8] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[7] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[6] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[5] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[4] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[3] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[2] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[1] = _zz_execute_ALUPlugin_subw_result;
    _zz_execute_ALUPlugin_subw_result_1[0] = _zz_execute_ALUPlugin_subw_result;
  end

  assign execute_ALUPlugin_subw_result = {_zz_execute_ALUPlugin_subw_result_1,_zz_execute_ALUPlugin_subw_result_2};
  assign execute_ALUPlugin_sllw_temp = (execute_ALUPlugin_src1_word <<< execute_ALUPlugin_shift_bits[4 : 0]);
  assign _zz_execute_ALUPlugin_sllw_result = execute_ALUPlugin_sllw_temp[31];
  always @(*) begin
    _zz_execute_ALUPlugin_sllw_result_1[31] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[30] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[29] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[28] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[27] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[26] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[25] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[24] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[23] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[22] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[21] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[20] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[19] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[18] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[17] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[16] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[15] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[14] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[13] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[12] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[11] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[10] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[9] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[8] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[7] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[6] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[5] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[4] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[3] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[2] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[1] = _zz_execute_ALUPlugin_sllw_result;
    _zz_execute_ALUPlugin_sllw_result_1[0] = _zz_execute_ALUPlugin_sllw_result;
  end

  assign execute_ALUPlugin_sllw_result = {_zz_execute_ALUPlugin_sllw_result_1,execute_ALUPlugin_sllw_temp};
  assign execute_ALUPlugin_srlw_temp = (execute_ALUPlugin_src1_word >>> execute_ALUPlugin_shift_bits[4 : 0]);
  assign _zz_execute_ALUPlugin_srlw_result = execute_ALUPlugin_srlw_temp[31];
  always @(*) begin
    _zz_execute_ALUPlugin_srlw_result_1[31] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[30] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[29] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[28] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[27] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[26] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[25] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[24] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[23] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[22] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[21] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[20] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[19] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[18] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[17] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[16] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[15] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[14] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[13] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[12] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[11] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[10] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[9] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[8] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[7] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[6] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[5] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[4] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[3] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[2] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[1] = _zz_execute_ALUPlugin_srlw_result;
    _zz_execute_ALUPlugin_srlw_result_1[0] = _zz_execute_ALUPlugin_srlw_result;
  end

  assign execute_ALUPlugin_srlw_result = {_zz_execute_ALUPlugin_srlw_result_1,execute_ALUPlugin_srlw_temp};
  assign execute_ALUPlugin_sraw_temp = ($signed(_zz_execute_ALUPlugin_sraw_temp) >>> execute_ALUPlugin_shift_bits[4 : 0]);
  assign _zz_execute_ALUPlugin_sraw_result = execute_ALUPlugin_sraw_temp[31];
  always @(*) begin
    _zz_execute_ALUPlugin_sraw_result_1[31] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[30] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[29] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[28] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[27] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[26] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[25] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[24] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[23] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[22] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[21] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[20] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[19] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[18] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[17] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[16] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[15] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[14] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[13] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[12] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[11] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[10] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[9] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[8] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[7] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[6] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[5] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[4] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[3] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[2] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[1] = _zz_execute_ALUPlugin_sraw_result;
    _zz_execute_ALUPlugin_sraw_result_1[0] = _zz_execute_ALUPlugin_sraw_result;
  end

  assign execute_ALUPlugin_sraw_result = {_zz_execute_ALUPlugin_sraw_result_1,execute_ALUPlugin_sraw_temp};
  assign execute_ALUPlugin_jal = (execute_ALU_CTRL == AluCtrlEnum_JAL);
  assign execute_ALUPlugin_jalr = (execute_ALU_CTRL == AluCtrlEnum_JALR);
  assign execute_ALUPlugin_beq = (execute_ALU_CTRL == AluCtrlEnum_BEQ);
  assign execute_ALUPlugin_bne = (execute_ALU_CTRL == AluCtrlEnum_BNE);
  assign execute_ALUPlugin_blt = (execute_ALU_CTRL == AluCtrlEnum_BLT);
  assign execute_ALUPlugin_bge = (execute_ALU_CTRL == AluCtrlEnum_BGE);
  assign execute_ALUPlugin_bltu = (execute_ALU_CTRL == AluCtrlEnum_BLTU);
  assign execute_ALUPlugin_bgeu = (execute_ALU_CTRL == AluCtrlEnum_BGEU);
  assign execute_ALUPlugin_branch_or_jalr = ((((((execute_ALUPlugin_jalr || execute_ALUPlugin_beq) || execute_ALUPlugin_bne) || execute_ALUPlugin_blt) || execute_ALUPlugin_bge) || execute_ALUPlugin_bltu) || execute_ALUPlugin_bgeu);
  assign execute_ALUPlugin_branch_or_jump = (execute_ALUPlugin_branch_or_jalr || execute_ALUPlugin_jal);
  assign execute_ALUPlugin_rd_is_link = ((execute_RD_ADDR == 5'h0) || (execute_RD_ADDR == 5'h05));
  assign execute_ALUPlugin_rs1_is_link = ((execute_RS1_ADDR == 5'h0) || (execute_RS1_ADDR == 5'h05));
  always @(*) begin
    execute_ALUPlugin_is_call = 1'b0;
    if(execute_ALUPlugin_jal) begin
      if(execute_ALUPlugin_rd_is_link) begin
        execute_ALUPlugin_is_call = 1'b1;
      end else begin
        execute_ALUPlugin_is_call = 1'b0;
      end
    end else begin
      if(execute_ALUPlugin_jalr) begin
        if(execute_ALUPlugin_rd_is_link) begin
          if(execute_ALUPlugin_rs1_is_link) begin
            if(when_AluPlugin_l270) begin
              execute_ALUPlugin_is_call = 1'b1;
            end else begin
              execute_ALUPlugin_is_call = 1'b1;
            end
          end else begin
            execute_ALUPlugin_is_call = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    execute_ALUPlugin_is_ret = 1'b0;
    if(execute_ALUPlugin_jal) begin
      if(execute_ALUPlugin_rd_is_link) begin
        execute_ALUPlugin_is_ret = 1'b0;
      end else begin
        execute_ALUPlugin_is_ret = 1'b0;
      end
    end else begin
      if(execute_ALUPlugin_jalr) begin
        if(execute_ALUPlugin_rd_is_link) begin
          if(execute_ALUPlugin_rs1_is_link) begin
            if(!when_AluPlugin_l270) begin
              execute_ALUPlugin_is_ret = 1'b1;
            end
          end
        end else begin
          if(execute_ALUPlugin_rs1_is_link) begin
            execute_ALUPlugin_is_ret = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    execute_ALUPlugin_is_jmp = 1'b0;
    if(execute_ALUPlugin_jal) begin
      if(execute_ALUPlugin_rd_is_link) begin
        execute_ALUPlugin_is_jmp = 1'b0;
      end else begin
        execute_ALUPlugin_is_jmp = 1'b1;
      end
    end else begin
      if(execute_ALUPlugin_jalr) begin
        if(!execute_ALUPlugin_rd_is_link) begin
          if(!execute_ALUPlugin_rs1_is_link) begin
            execute_ALUPlugin_is_jmp = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    execute_ALUPlugin_redirect_pc_next = (execute_PC + 64'h0000000000000004);
    if(execute_ALUPlugin_branch_or_jump) begin
      if(execute_ALUPlugin_branch_taken) begin
        if(when_AluPlugin_l234) begin
          execute_ALUPlugin_redirect_pc_next = execute_ALUPlugin_pc_next;
        end
      end else begin
        if(execute_PREDICT_TAKEN) begin
          execute_ALUPlugin_redirect_pc_next = (execute_PC + 64'h0000000000000004);
        end
      end
    end
  end

  always @(*) begin
    execute_ALUPlugin_redirect_valid = 1'b0;
    if(execute_ALUPlugin_branch_or_jump) begin
      if(execute_ALUPlugin_branch_taken) begin
        if(when_AluPlugin_l234) begin
          execute_ALUPlugin_redirect_valid = execute_arbitration_isFiring;
        end
      end else begin
        if(execute_PREDICT_TAKEN) begin
          execute_ALUPlugin_redirect_valid = execute_arbitration_isFiring;
        end
      end
    end
  end

  assign when_AluPlugin_l77 = (((execute_ALU_CTRL == AluCtrlEnum_AUIPC) || execute_ALUPlugin_jal) || execute_ALUPlugin_jalr);
  always @(*) begin
    if(when_AluPlugin_l77) begin
      execute_ALUPlugin_src1 = execute_PC;
    end else begin
      if(execute_RS1_FROM_MEM) begin
        execute_ALUPlugin_src1 = memaccess_ALU_RESULT;
      end else begin
        if(execute_RS1_FROM_LOAD) begin
          execute_ALUPlugin_src1 = memaccess_LSU_RDATA;
        end else begin
          if(execute_RS1_FROM_WB) begin
            execute_ALUPlugin_src1 = _zz_execute_MEM_WDATA_2;
          end else begin
            execute_ALUPlugin_src1 = execute_RS1;
          end
        end
      end
    end
  end

  assign when_AluPlugin_l95 = (execute_ALUPlugin_jal || execute_ALUPlugin_jalr);
  always @(*) begin
    if(when_AluPlugin_l95) begin
      execute_ALUPlugin_src2 = 64'h0000000000000004;
    end else begin
      if(execute_SRC2_IS_IMM) begin
        execute_ALUPlugin_src2 = execute_IMM;
      end else begin
        if(execute_RS2_FROM_MEM) begin
          execute_ALUPlugin_src2 = memaccess_ALU_RESULT;
        end else begin
          if(execute_RS2_FROM_LOAD) begin
            execute_ALUPlugin_src2 = memaccess_LSU_RDATA;
          end else begin
            if(execute_RS2_FROM_WB) begin
              execute_ALUPlugin_src2 = _zz_execute_MEM_WDATA_2;
            end else begin
              execute_ALUPlugin_src2 = execute_RS2;
            end
          end
        end
      end
    end
  end

  always @(*) begin
    if(execute_CTRL_RS1_FROM_MEM) begin
      execute_ALUPlugin_branch_src1 = _zz_execute_MEM_WDATA_1;
    end else begin
      if(execute_CTRL_RS1_FROM_LOAD) begin
        execute_ALUPlugin_branch_src1 = _zz_execute_MEM_WDATA;
      end else begin
        if(execute_CTRL_RS1_FROM_WB) begin
          execute_ALUPlugin_branch_src1 = _zz_execute_MEM_WDATA_2;
        end else begin
          execute_ALUPlugin_branch_src1 = execute_RS1;
        end
      end
    end
  end

  always @(*) begin
    if(execute_CTRL_RS2_FROM_MEM) begin
      execute_ALUPlugin_branch_src2 = _zz_execute_MEM_WDATA_1;
    end else begin
      if(execute_CTRL_RS2_FROM_LOAD) begin
        execute_ALUPlugin_branch_src2 = _zz_execute_MEM_WDATA;
      end else begin
        if(execute_CTRL_RS2_FROM_WB) begin
          execute_ALUPlugin_branch_src2 = _zz_execute_MEM_WDATA_2;
        end else begin
          execute_ALUPlugin_branch_src2 = execute_RS2;
        end
      end
    end
  end

  assign when_AluPlugin_l146 = (execute_ALU_WORD == 1'b1);
  always @(*) begin
    if((execute_ALU_CTRL == AluCtrlEnum_ADD)) begin
        if(when_AluPlugin_l146) begin
          execute_ALUPlugin_alu_result = execute_ALUPlugin_addw_result;
        end else begin
          execute_ALUPlugin_alu_result = execute_ALUPlugin_add_result;
        end
    end else if((execute_ALU_CTRL == AluCtrlEnum_SUB)) begin
        if(when_AluPlugin_l153) begin
          execute_ALUPlugin_alu_result = execute_ALUPlugin_subw_result;
        end else begin
          execute_ALUPlugin_alu_result = execute_ALUPlugin_sub_result;
        end
    end else if((execute_ALU_CTRL == AluCtrlEnum_SLT)) begin
        execute_ALUPlugin_alu_result = {_zz_execute_ALUPlugin_alu_result,execute_ALUPlugin_slt_result};
    end else if((execute_ALU_CTRL == AluCtrlEnum_SLTU)) begin
        execute_ALUPlugin_alu_result = {_zz_execute_ALUPlugin_alu_result_1,execute_ALUPlugin_sltu_result};
    end else if((execute_ALU_CTRL == AluCtrlEnum_XOR_1)) begin
        execute_ALUPlugin_alu_result = execute_ALUPlugin_xor_result;
    end else if((execute_ALU_CTRL == AluCtrlEnum_SLL_1)) begin
        if(when_AluPlugin_l169) begin
          execute_ALUPlugin_alu_result = execute_ALUPlugin_sllw_result;
        end else begin
          execute_ALUPlugin_alu_result = execute_ALUPlugin_sll_result;
        end
    end else if((execute_ALU_CTRL == AluCtrlEnum_SRL_1)) begin
        if(when_AluPlugin_l176) begin
          execute_ALUPlugin_alu_result = execute_ALUPlugin_srlw_result;
        end else begin
          execute_ALUPlugin_alu_result = execute_ALUPlugin_srl_result;
        end
    end else if((execute_ALU_CTRL == AluCtrlEnum_SRA_1)) begin
        if(when_AluPlugin_l183) begin
          execute_ALUPlugin_alu_result = execute_ALUPlugin_sraw_result;
        end else begin
          execute_ALUPlugin_alu_result = execute_ALUPlugin_sra_result;
        end
    end else if((execute_ALU_CTRL == AluCtrlEnum_AND_1)) begin
        execute_ALUPlugin_alu_result = execute_ALUPlugin_and_result;
    end else if((execute_ALU_CTRL == AluCtrlEnum_OR_1)) begin
        execute_ALUPlugin_alu_result = execute_ALUPlugin_or_result;
    end else if((execute_ALU_CTRL == AluCtrlEnum_LUI)) begin
        execute_ALUPlugin_alu_result = execute_IMM;
    end else if((execute_ALU_CTRL == AluCtrlEnum_JAL) || (execute_ALU_CTRL == AluCtrlEnum_JALR) || (execute_ALU_CTRL == AluCtrlEnum_AUIPC)) begin
        execute_ALUPlugin_alu_result = execute_ALUPlugin_add_result;
    end else if((execute_ALU_CTRL == AluCtrlEnum_CSR)) begin
        execute_ALUPlugin_alu_result = execute_CSR_RDATA;
    end else begin
        execute_ALUPlugin_alu_result = execute_ALUPlugin_add_result;
    end
  end

  assign when_AluPlugin_l153 = (execute_ALU_WORD == 1'b1);
  assign _zz_execute_ALUPlugin_alu_result[62 : 0] = 63'h0;
  assign _zz_execute_ALUPlugin_alu_result_1[62 : 0] = 63'h0;
  assign when_AluPlugin_l169 = (execute_ALU_WORD == 1'b1);
  assign when_AluPlugin_l176 = (execute_ALU_WORD == 1'b1);
  assign when_AluPlugin_l183 = (execute_ALU_WORD == 1'b1);
  assign execute_ALUPlugin_beq_result = (execute_ALUPlugin_beq && (execute_ALUPlugin_branch_src1 == execute_ALUPlugin_branch_src2));
  assign execute_ALUPlugin_bne_result = (execute_ALUPlugin_bne && (execute_ALUPlugin_branch_src1 != execute_ALUPlugin_branch_src2));
  assign execute_ALUPlugin_blt_result = (execute_ALUPlugin_blt && ($signed(_zz_execute_ALUPlugin_blt_result) < $signed(_zz_execute_ALUPlugin_blt_result_1)));
  assign execute_ALUPlugin_bge_result = (execute_ALUPlugin_bge && ($signed(_zz_execute_ALUPlugin_bge_result) <= $signed(_zz_execute_ALUPlugin_bge_result_1)));
  assign execute_ALUPlugin_bltu_result = (execute_ALUPlugin_bltu && (execute_ALUPlugin_branch_src1 < execute_ALUPlugin_branch_src2));
  assign execute_ALUPlugin_bgeu_result = (execute_ALUPlugin_bgeu && (execute_ALUPlugin_branch_src2 <= execute_ALUPlugin_branch_src1));
  assign execute_ALUPlugin_branch_taken = (((((((execute_ALUPlugin_beq_result || execute_ALUPlugin_bne_result) || execute_ALUPlugin_blt_result) || execute_ALUPlugin_bge_result) || execute_ALUPlugin_bltu_result) || execute_ALUPlugin_bgeu_result) || execute_ALUPlugin_jal) || execute_ALUPlugin_jalr);
  assign when_AluPlugin_l226 = (execute_ALU_CTRL == AluCtrlEnum_JALR);
  always @(*) begin
    if(when_AluPlugin_l226) begin
      execute_ALUPlugin_pc_next = _zz_execute_ALUPlugin_pc_next;
    end else begin
      execute_ALUPlugin_pc_next = _zz_execute_ALUPlugin_pc_next_6;
    end
  end

  assign when_AluPlugin_l234 = ((! execute_PREDICT_TAKEN) || (execute_PC_NEXT != execute_ALUPlugin_pc_next));
  assign when_AluPlugin_l270 = (execute_RD_ADDR == execute_RS1_ADDR);
  assign DecodePlugin_hazard_rs1_from_mem = ((((memaccess_arbitration_isValid && _zz_DecodePlugin_hazard_rs1_from_mem_3) && (_zz_DecodePlugin_hazard_rs1_from_mem_2 != 5'h0)) && (_zz_DecodePlugin_hazard_rs1_from_mem_2 == _zz_DecodePlugin_hazard_rs1_from_mem_1)) && (! _zz_DecodePlugin_hazard_rs1_from_mem));
  assign DecodePlugin_hazard_rs2_from_mem = ((((memaccess_arbitration_isValid && _zz_DecodePlugin_hazard_rs1_from_mem_3) && (_zz_DecodePlugin_hazard_rs1_from_mem_2 != 5'h0)) && (_zz_DecodePlugin_hazard_rs1_from_mem_2 == _zz_DecodePlugin_hazard_rs2_from_mem)) && (! _zz_DecodePlugin_hazard_rs1_from_mem));
  assign DecodePlugin_hazard_rs1_from_load = ((((memaccess_arbitration_isValid && _zz_DecodePlugin_hazard_rs1_from_mem_3) && (_zz_DecodePlugin_hazard_rs1_from_mem_2 != 5'h0)) && (_zz_DecodePlugin_hazard_rs1_from_mem_2 == _zz_DecodePlugin_hazard_rs1_from_mem_1)) && _zz_DecodePlugin_hazard_rs1_from_mem);
  assign DecodePlugin_hazard_rs2_from_load = ((((memaccess_arbitration_isValid && _zz_DecodePlugin_hazard_rs1_from_mem_3) && (_zz_DecodePlugin_hazard_rs1_from_mem_2 != 5'h0)) && (_zz_DecodePlugin_hazard_rs1_from_mem_2 == _zz_DecodePlugin_hazard_rs2_from_mem)) && _zz_DecodePlugin_hazard_rs1_from_mem);
  assign DecodePlugin_hazard_rs1_from_wb = ((((writeback_arbitration_isValid && _zz_DecodePlugin_hazard_rs1_from_wb_1) && (_zz_DecodePlugin_hazard_rs1_from_wb != 5'h0)) && (_zz_DecodePlugin_hazard_rs1_from_wb == _zz_DecodePlugin_hazard_rs1_from_mem_1)) && (! (DecodePlugin_hazard_rs1_from_mem || DecodePlugin_hazard_rs1_from_load)));
  assign DecodePlugin_hazard_rs2_from_wb = ((((writeback_arbitration_isValid && _zz_DecodePlugin_hazard_rs1_from_wb_1) && (_zz_DecodePlugin_hazard_rs1_from_wb != 5'h0)) && (_zz_DecodePlugin_hazard_rs1_from_wb == _zz_DecodePlugin_hazard_rs2_from_mem)) && (! (DecodePlugin_hazard_rs2_from_mem || DecodePlugin_hazard_rs2_from_load)));
  assign DecodePlugin_hazard_load_use = ((memaccess_arbitration_isValid && _zz_DecodePlugin_hazard_rs1_from_mem) && (((_zz_DecodePlugin_hazard_rs1_from_mem_2 == _zz_DecodePlugin_hazard_rs1_from_mem_1) && (! DecodePlugin_hazard_rs1_from_wb)) || ((_zz_DecodePlugin_hazard_rs1_from_mem_2 == _zz_DecodePlugin_hazard_rs2_from_mem) && (! DecodePlugin_hazard_rs2_from_wb))));
  assign DecodePlugin_hazard_ctrl_rs1_from_mem = ((execute_arbitration_isValid && _zz_DecodePlugin_hazard_ctrl_rs1_from_mem) && DecodePlugin_hazard_rs1_from_mem);
  assign DecodePlugin_hazard_ctrl_rs2_from_mem = ((execute_arbitration_isValid && _zz_DecodePlugin_hazard_ctrl_rs1_from_mem) && DecodePlugin_hazard_rs2_from_mem);
  assign DecodePlugin_hazard_ctrl_rs1_from_load = ((execute_arbitration_isValid && _zz_DecodePlugin_hazard_ctrl_rs1_from_mem) && DecodePlugin_hazard_rs1_from_load);
  assign DecodePlugin_hazard_ctrl_rs2_from_load = ((execute_arbitration_isValid && _zz_DecodePlugin_hazard_ctrl_rs1_from_mem) && DecodePlugin_hazard_rs2_from_load);
  assign DecodePlugin_hazard_ctrl_rs1_from_wb = ((execute_arbitration_isValid && _zz_DecodePlugin_hazard_ctrl_rs1_from_mem) && DecodePlugin_hazard_rs1_from_wb);
  assign DecodePlugin_hazard_ctrl_rs2_from_wb = ((execute_arbitration_isValid && _zz_DecodePlugin_hazard_ctrl_rs1_from_mem) && DecodePlugin_hazard_rs2_from_wb);
  assign DecodePlugin_hazard_ctrl_load_use = ((execute_arbitration_isValid && _zz_DecodePlugin_hazard_ctrl_rs1_from_mem) && DecodePlugin_hazard_load_use);
  assign fetch_arbitration_haltItself = 1'b0;
  assign fetch_arbitration_flushIt = (when_FetchPlugin_l97 || when_FetchPlugin_l94);
  assign decode_arbitration_haltItself = 1'b0;
  assign decode_arbitration_flushIt = (when_FetchPlugin_l97 || when_FetchPlugin_l94);
  assign execute_arbitration_haltItself = execute_INT_HOLD;
  assign execute_arbitration_flushIt = 1'b0;
  assign memaccess_arbitration_haltItself = _zz_memaccess_arbitration_haltItself;
  assign memaccess_arbitration_flushIt = 1'b0;
  assign writeback_arbitration_haltItself = _zz_memaccess_arbitration_haltItself;
  assign writeback_arbitration_flushIt = 1'b0;
  assign clint_1_ecall = (execute_arbitration_isValid && (_zz_ecall == CsrCtrlEnum_ECALL));
  assign clint_1_ebreak = (execute_arbitration_isValid && (_zz_ecall == CsrCtrlEnum_EBREAK));
  assign clint_1_mret = (execute_arbitration_isValid && (_zz_ecall == CsrCtrlEnum_MRET));
  assign execute_ExcepPlugin_csrrs_wdata = (execute_SRC1 | execute_CSR_RDATA);
  assign execute_ExcepPlugin_csrrc_wdata = ((~ execute_SRC1) & execute_CSR_RDATA);
  assign execute_ExcepPlugin_csrrsi_wdata = (execute_IMM | execute_CSR_RDATA);
  assign execute_ExcepPlugin_csrrci_wdata = ((~ execute_IMM) & execute_CSR_RDATA);
  always @(*) begin
    if((execute_CSR_CTRL == CsrCtrlEnum_CSRRW)) begin
        execute_ExcepPlugin_csr_wdata = execute_SRC1;
    end else if((execute_CSR_CTRL == CsrCtrlEnum_CSRRS)) begin
        execute_ExcepPlugin_csr_wdata = execute_ExcepPlugin_csrrs_wdata;
    end else if((execute_CSR_CTRL == CsrCtrlEnum_CSRRC)) begin
        execute_ExcepPlugin_csr_wdata = execute_ExcepPlugin_csrrc_wdata;
    end else if((execute_CSR_CTRL == CsrCtrlEnum_CSRRWI)) begin
        execute_ExcepPlugin_csr_wdata = execute_IMM;
    end else if((execute_CSR_CTRL == CsrCtrlEnum_CSRRSI)) begin
        execute_ExcepPlugin_csr_wdata = execute_ExcepPlugin_csrrsi_wdata;
    end else if((execute_CSR_CTRL == CsrCtrlEnum_CSRRCI)) begin
        execute_ExcepPlugin_csr_wdata = execute_ExcepPlugin_csrrci_wdata;
    end else begin
        execute_ExcepPlugin_csr_wdata = 64'h0;
    end
  end

  assign timer_1_addr = _zz_execute_MEM_WDATA_1;
  assign memaccess_LSUPlugin_cpu_addr = memaccess_ALU_RESULT;
  assign memaccess_LSUPlugin_cpu_addr_offset = memaccess_LSUPlugin_cpu_addr[2 : 0];
  assign memaccess_LSUPlugin_is_mem = (memaccess_IS_LOAD || memaccess_IS_STORE);
  assign memaccess_LSUPlugin_is_timer = ((memaccess_LSUPlugin_cpu_addr == 64'h000000000200bff8) || (memaccess_LSUPlugin_cpu_addr == 64'h0000000002004000));
  assign memaccess_LSUPlugin_dcache_rdata = (DCachePlugin_dcache_access_rsp_payload_data >>> _zz_memaccess_LSUPlugin_dcache_rdata);
  assign _zz_memaccess_LSUPlugin_dcache_lb = memaccess_LSUPlugin_dcache_rdata[7];
  always @(*) begin
    _zz_memaccess_LSUPlugin_dcache_lb_1[55] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[54] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[53] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[52] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[51] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[50] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[49] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[48] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[47] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[46] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[45] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[44] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[43] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[42] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[41] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[40] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[39] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[38] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[37] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[36] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[35] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[34] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[33] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[32] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[31] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[30] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[29] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[28] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[27] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[26] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[25] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[24] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[23] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[22] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[21] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[20] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[19] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[18] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[17] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[16] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[15] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[14] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[13] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[12] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[11] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[10] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[9] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[8] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[7] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[6] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[5] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[4] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[3] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[2] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[1] = _zz_memaccess_LSUPlugin_dcache_lb;
    _zz_memaccess_LSUPlugin_dcache_lb_1[0] = _zz_memaccess_LSUPlugin_dcache_lb;
  end

  assign memaccess_LSUPlugin_dcache_lb = {_zz_memaccess_LSUPlugin_dcache_lb_1,memaccess_LSUPlugin_dcache_rdata[7 : 0]};
  assign _zz_1 = zz__zz_memaccess_LSUPlugin_dcache_lbu(1'b0);
  always @(*) _zz_memaccess_LSUPlugin_dcache_lbu = _zz_1;
  assign memaccess_LSUPlugin_dcache_lbu = {_zz_memaccess_LSUPlugin_dcache_lbu,memaccess_LSUPlugin_dcache_rdata[7 : 0]};
  assign _zz_memaccess_LSUPlugin_dcache_lh = memaccess_LSUPlugin_dcache_rdata[15];
  always @(*) begin
    _zz_memaccess_LSUPlugin_dcache_lh_1[47] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[46] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[45] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[44] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[43] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[42] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[41] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[40] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[39] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[38] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[37] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[36] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[35] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[34] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[33] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[32] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[31] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[30] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[29] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[28] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[27] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[26] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[25] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[24] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[23] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[22] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[21] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[20] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[19] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[18] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[17] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[16] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[15] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[14] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[13] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[12] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[11] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[10] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[9] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[8] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[7] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[6] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[5] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[4] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[3] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[2] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[1] = _zz_memaccess_LSUPlugin_dcache_lh;
    _zz_memaccess_LSUPlugin_dcache_lh_1[0] = _zz_memaccess_LSUPlugin_dcache_lh;
  end

  assign memaccess_LSUPlugin_dcache_lh = {_zz_memaccess_LSUPlugin_dcache_lh_1,memaccess_LSUPlugin_dcache_rdata[15 : 0]};
  assign _zz_2 = zz__zz_memaccess_LSUPlugin_dcache_lhu(1'b0);
  always @(*) _zz_memaccess_LSUPlugin_dcache_lhu = _zz_2;
  assign memaccess_LSUPlugin_dcache_lhu = {_zz_memaccess_LSUPlugin_dcache_lhu,memaccess_LSUPlugin_dcache_rdata[15 : 0]};
  assign _zz_memaccess_LSUPlugin_dcache_lw = memaccess_LSUPlugin_dcache_rdata[31];
  always @(*) begin
    _zz_memaccess_LSUPlugin_dcache_lw_1[31] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[30] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[29] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[28] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[27] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[26] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[25] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[24] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[23] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[22] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[21] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[20] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[19] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[18] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[17] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[16] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[15] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[14] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[13] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[12] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[11] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[10] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[9] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[8] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[7] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[6] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[5] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[4] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[3] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[2] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[1] = _zz_memaccess_LSUPlugin_dcache_lw;
    _zz_memaccess_LSUPlugin_dcache_lw_1[0] = _zz_memaccess_LSUPlugin_dcache_lw;
  end

  assign memaccess_LSUPlugin_dcache_lw = {_zz_memaccess_LSUPlugin_dcache_lw_1,memaccess_LSUPlugin_dcache_rdata[31 : 0]};
  assign _zz_3 = zz__zz_memaccess_LSUPlugin_dcache_lwu(1'b0);
  always @(*) _zz_memaccess_LSUPlugin_dcache_lwu = _zz_3;
  assign memaccess_LSUPlugin_dcache_lwu = {_zz_memaccess_LSUPlugin_dcache_lwu,memaccess_LSUPlugin_dcache_rdata[31 : 0]};
  assign _zz_memaccess_LSUPlugin_dcache_sb = memaccess_MEM_WDATA[7];
  always @(*) begin
    _zz_memaccess_LSUPlugin_dcache_sb_1[55] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[54] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[53] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[52] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[51] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[50] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[49] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[48] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[47] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[46] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[45] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[44] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[43] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[42] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[41] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[40] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[39] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[38] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[37] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[36] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[35] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[34] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[33] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[32] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[31] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[30] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[29] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[28] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[27] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[26] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[25] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[24] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[23] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[22] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[21] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[20] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[19] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[18] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[17] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[16] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[15] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[14] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[13] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[12] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[11] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[10] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[9] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[8] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[7] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[6] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[5] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[4] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[3] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[2] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[1] = _zz_memaccess_LSUPlugin_dcache_sb;
    _zz_memaccess_LSUPlugin_dcache_sb_1[0] = _zz_memaccess_LSUPlugin_dcache_sb;
  end

  assign memaccess_LSUPlugin_dcache_sb = {_zz_memaccess_LSUPlugin_dcache_sb_1,memaccess_MEM_WDATA[7 : 0]};
  assign _zz_memaccess_LSUPlugin_dcache_sh = memaccess_MEM_WDATA[15];
  always @(*) begin
    _zz_memaccess_LSUPlugin_dcache_sh_1[47] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[46] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[45] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[44] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[43] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[42] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[41] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[40] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[39] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[38] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[37] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[36] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[35] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[34] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[33] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[32] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[31] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[30] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[29] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[28] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[27] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[26] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[25] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[24] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[23] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[22] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[21] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[20] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[19] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[18] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[17] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[16] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[15] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[14] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[13] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[12] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[11] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[10] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[9] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[8] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[7] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[6] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[5] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[4] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[3] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[2] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[1] = _zz_memaccess_LSUPlugin_dcache_sh;
    _zz_memaccess_LSUPlugin_dcache_sh_1[0] = _zz_memaccess_LSUPlugin_dcache_sh;
  end

  assign memaccess_LSUPlugin_dcache_sh = {_zz_memaccess_LSUPlugin_dcache_sh_1,memaccess_MEM_WDATA[15 : 0]};
  assign _zz_memaccess_LSUPlugin_dcache_sw = memaccess_MEM_WDATA[31];
  always @(*) begin
    _zz_memaccess_LSUPlugin_dcache_sw_1[31] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[30] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[29] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[28] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[27] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[26] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[25] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[24] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[23] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[22] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[21] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[20] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[19] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[18] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[17] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[16] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[15] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[14] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[13] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[12] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[11] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[10] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[9] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[8] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[7] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[6] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[5] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[4] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[3] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[2] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[1] = _zz_memaccess_LSUPlugin_dcache_sw;
    _zz_memaccess_LSUPlugin_dcache_sw_1[0] = _zz_memaccess_LSUPlugin_dcache_sw;
  end

  assign memaccess_LSUPlugin_dcache_sw = {_zz_memaccess_LSUPlugin_dcache_sw_1,memaccess_MEM_WDATA[31 : 0]};
  assign memaccess_LSUPlugin_lsu_ready = 1'b1;
  always @(*) begin
    if((memaccess_MEM_CTRL == MemCtrlEnum_LB)) begin
        memaccess_LSUPlugin_dcache_data_load = memaccess_LSUPlugin_dcache_lb;
    end else if((memaccess_MEM_CTRL == MemCtrlEnum_LBU)) begin
        memaccess_LSUPlugin_dcache_data_load = memaccess_LSUPlugin_dcache_lbu;
    end else if((memaccess_MEM_CTRL == MemCtrlEnum_LH)) begin
        memaccess_LSUPlugin_dcache_data_load = memaccess_LSUPlugin_dcache_lh;
    end else if((memaccess_MEM_CTRL == MemCtrlEnum_LHU)) begin
        memaccess_LSUPlugin_dcache_data_load = memaccess_LSUPlugin_dcache_lhu;
    end else if((memaccess_MEM_CTRL == MemCtrlEnum_LW)) begin
        memaccess_LSUPlugin_dcache_data_load = memaccess_LSUPlugin_dcache_lw;
    end else if((memaccess_MEM_CTRL == MemCtrlEnum_LWU)) begin
        memaccess_LSUPlugin_dcache_data_load = memaccess_LSUPlugin_dcache_lwu;
    end else if((memaccess_MEM_CTRL == MemCtrlEnum_LD)) begin
        memaccess_LSUPlugin_dcache_data_load = memaccess_LSUPlugin_dcache_rdata;
    end else begin
        memaccess_LSUPlugin_dcache_data_load = 64'h0;
    end
  end

  always @(*) begin
    if((memaccess_MEM_CTRL == MemCtrlEnum_SB)) begin
        memaccess_LSUPlugin_dcache_wdata = memaccess_LSUPlugin_dcache_sb;
    end else if((memaccess_MEM_CTRL == MemCtrlEnum_SH)) begin
        memaccess_LSUPlugin_dcache_wdata = memaccess_LSUPlugin_dcache_sh;
    end else if((memaccess_MEM_CTRL == MemCtrlEnum_SW)) begin
        memaccess_LSUPlugin_dcache_wdata = memaccess_LSUPlugin_dcache_sw;
    end else if((memaccess_MEM_CTRL == MemCtrlEnum_SD)) begin
        memaccess_LSUPlugin_dcache_wdata = memaccess_MEM_WDATA;
    end else begin
        memaccess_LSUPlugin_dcache_wdata = 64'h0;
    end
  end

  assign _zz_4 = zz__zz_memaccess_LSUPlugin_dcache_wstrb(1'b0);
  always @(*) _zz_memaccess_LSUPlugin_dcache_wstrb = _zz_4;
  always @(*) begin
    if((memaccess_MEM_CTRL == MemCtrlEnum_SB)) begin
        memaccess_LSUPlugin_dcache_wstrb = _zz_memaccess_LSUPlugin_dcache_wstrb;
    end else if((memaccess_MEM_CTRL == MemCtrlEnum_SH)) begin
        memaccess_LSUPlugin_dcache_wstrb = _zz_memaccess_LSUPlugin_dcache_wstrb_1;
    end else if((memaccess_MEM_CTRL == MemCtrlEnum_SW)) begin
        memaccess_LSUPlugin_dcache_wstrb = _zz_memaccess_LSUPlugin_dcache_wstrb_2;
    end else if((memaccess_MEM_CTRL == MemCtrlEnum_SD)) begin
        memaccess_LSUPlugin_dcache_wstrb = _zz_memaccess_LSUPlugin_dcache_wstrb_3;
    end else begin
        memaccess_LSUPlugin_dcache_wstrb = 8'h0;
    end
  end

  assign _zz_5 = zz__zz_memaccess_LSUPlugin_dcache_wstrb_1(1'b0);
  always @(*) _zz_memaccess_LSUPlugin_dcache_wstrb_1 = _zz_5;
  assign _zz_6 = zz__zz_memaccess_LSUPlugin_dcache_wstrb_2(1'b0);
  always @(*) _zz_memaccess_LSUPlugin_dcache_wstrb_2 = _zz_6;
  assign _zz_memaccess_LSUPlugin_dcache_wstrb_3[7 : 0] = 8'hff;
  assign memaccess_LSUPlugin_lsu_rdata = memaccess_LSUPlugin_dcache_data_load;
  assign memaccess_LSUPlugin_lsu_wdata = (memaccess_LSUPlugin_dcache_wdata <<< _zz_memaccess_LSUPlugin_lsu_wdata);
  assign memaccess_LSUPlugin_lsu_addr = memaccess_LSUPlugin_cpu_addr;
  assign memaccess_LSUPlugin_lsu_wen = memaccess_IS_STORE;
  assign memaccess_LSUPlugin_lsu_wstrb = (memaccess_LSUPlugin_dcache_wstrb <<< memaccess_LSUPlugin_cpu_addr_offset);
  assign DCachePlugin_dcache_access_cmd_valid = (((! memaccess_LSUPlugin_is_timer) && memaccess_LSUPlugin_is_mem) && memaccess_arbitration_isValid);
  assign DCachePlugin_dcache_access_cmd_payload_addr = memaccess_LSUPlugin_lsu_addr;
  assign DCachePlugin_dcache_access_cmd_payload_wen = memaccess_LSUPlugin_lsu_wen;
  assign DCachePlugin_dcache_access_cmd_payload_wdata = memaccess_LSUPlugin_lsu_wdata;
  assign DCachePlugin_dcache_access_cmd_payload_wstrb = memaccess_LSUPlugin_lsu_wstrb;
  assign ICachePlugin_icache_access_cmd_ready = iCache_1_cpu_cmd_ready;
  assign ICachePlugin_icache_access_rsp_valid = iCache_1_cpu_rsp_valid;
  assign ICachePlugin_icache_access_rsp_payload_data = iCache_1_cpu_rsp_payload_data;
  assign icache_ar_valid = iCache_1_next_level_cmd_valid;
  assign icache_ar_payload_id = 4'b0000;
  assign icache_ar_payload_len = {4'd0, iCache_1_next_level_cmd_payload_len};
  assign icache_ar_payload_size = iCache_1_next_level_cmd_payload_size;
  assign icache_ar_payload_burst = 2'b01;
  assign icache_ar_payload_addr = iCache_1_next_level_cmd_payload_addr;
  assign icache_r_ready = 1'b1;
  assign DCachePlugin_dcache_access_cmd_ready = dCache_1_cpu_cmd_ready;
  assign DCachePlugin_dcache_access_rsp_valid = dCache_1_cpu_rsp_valid;
  assign DCachePlugin_dcache_access_rsp_payload_data = dCache_1_cpu_rsp_payload_data;
  assign DCachePlugin_dcache_access_stall = dCache_1_stall;
  assign when_DCachePlugin_l118 = (dCache_1_next_level_cmd_valid && (! dCache_1_next_level_cmd_payload_wen));
  assign dcache_ar_fire = (dcache_ar_valid && dcache_ar_ready);
  assign dcache_r_ready = 1'b1;
  assign when_DCachePlugin_l141 = (dCache_1_next_level_cmd_valid && dCache_1_next_level_cmd_payload_wen);
  assign dcache_aw_fire = (dcache_aw_valid && dcache_aw_ready);
  assign when_DCachePlugin_l159 = (dCache_1_next_level_cmd_valid && dCache_1_next_level_cmd_payload_wen);
  assign dcache_w_fire = (dcache_w_valid && dcache_w_ready);
  assign dcache_b_ready = 1'b1;
  assign when_DCachePlugin_l174 = (_zz_when_DCachePlugin_l174 == 1'b0);
  assign dcache_aw_fire_1 = (dcache_aw_valid && dcache_aw_ready);
  assign dcache_w_fire_1 = (dcache_w_valid && dcache_w_ready);
  assign when_DCachePlugin_l175 = (dcache_aw_fire_1 && dcache_w_fire_1);
  assign dcache_aw_fire_2 = (dcache_aw_valid && dcache_aw_ready);
  assign dcache_w_fire_2 = (dcache_w_valid && dcache_w_ready);
  assign when_DCachePlugin_l177 = (dcache_aw_fire_2 || dcache_w_fire_2);
  assign dcache_aw_fire_3 = (dcache_aw_valid && dcache_aw_ready);
  assign dcache_w_fire_3 = (dcache_w_valid && dcache_w_ready);
  assign when_DCachePlugin_l182 = (dcache_aw_fire_3 || dcache_w_fire_3);
  assign when_DCachePlugin_l181 = (_zz_when_DCachePlugin_l174 == 1'b1);
  assign dcache_aw_fire_4 = (dcache_aw_valid && dcache_aw_ready);
  assign dcache_w_fire_4 = (dcache_w_valid && dcache_w_ready);
  assign dcache_aw_fire_5 = (dcache_aw_valid && dcache_aw_ready);
  assign dcache_w_fire_5 = (dcache_w_valid && dcache_w_ready);
  assign dCache_1_next_level_cmd_ready = (dCache_1_next_level_cmd_payload_wen ? ((dcache_aw_fire_4 && dcache_w_fire_4) || (_zz_when_DCachePlugin_l174 && (dcache_aw_fire_5 || dcache_w_fire_5))) : dcache_ar_ready);
  assign dCache_1_next_level_rsp_valid = (dCache_1_next_level_cmd_payload_wen ? dcache_b_valid : dcache_r_valid);
  assign when_Pipeline_l127 = (! decode_arbitration_isStuck);
  assign when_Pipeline_l127_1 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_2 = (! memaccess_arbitration_isStuck);
  assign when_Pipeline_l127_3 = (! writeback_arbitration_isStuck);
  assign when_Pipeline_l127_4 = (! decode_arbitration_isStuck);
  assign when_Pipeline_l127_5 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_6 = (! decode_arbitration_isStuck);
  assign when_Pipeline_l127_7 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_8 = (! memaccess_arbitration_isStuck);
  assign when_Pipeline_l127_9 = (! writeback_arbitration_isStuck);
  assign when_Pipeline_l127_10 = (! decode_arbitration_isStuck);
  assign when_Pipeline_l127_11 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_12 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_13 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_14 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_15 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_16 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_17 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_18 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_19 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_20 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_21 = (! memaccess_arbitration_isStuck);
  assign when_Pipeline_l127_22 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_23 = (! memaccess_arbitration_isStuck);
  assign when_Pipeline_l127_24 = (! writeback_arbitration_isStuck);
  assign when_Pipeline_l127_25 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_26 = (! memaccess_arbitration_isStuck);
  assign when_Pipeline_l127_27 = (! writeback_arbitration_isStuck);
  assign when_Pipeline_l127_28 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_29 = (! memaccess_arbitration_isStuck);
  assign when_Pipeline_l127_30 = (! writeback_arbitration_isStuck);
  assign when_Pipeline_l127_31 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_32 = (! memaccess_arbitration_isStuck);
  assign when_Pipeline_l127_33 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_34 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_35 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_36 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l127_37 = (! memaccess_arbitration_isStuck);
  assign when_Pipeline_l127_38 = (! writeback_arbitration_isStuck);
  assign when_Pipeline_l127_39 = (! memaccess_arbitration_isStuck);
  assign when_Pipeline_l127_40 = (! writeback_arbitration_isStuck);
  assign fetch_arbitration_isFlushed = (({writeback_arbitration_flushNext,{memaccess_arbitration_flushNext,{execute_arbitration_flushNext,decode_arbitration_flushNext}}} != 4'b0000) || ({writeback_arbitration_flushIt,{memaccess_arbitration_flushIt,{execute_arbitration_flushIt,{decode_arbitration_flushIt,fetch_arbitration_flushIt}}}} != 5'h0));
  assign decode_arbitration_isFlushed = (({writeback_arbitration_flushNext,{memaccess_arbitration_flushNext,execute_arbitration_flushNext}} != 3'b000) || ({writeback_arbitration_flushIt,{memaccess_arbitration_flushIt,{execute_arbitration_flushIt,decode_arbitration_flushIt}}} != 4'b0000));
  assign execute_arbitration_isFlushed = (({writeback_arbitration_flushNext,memaccess_arbitration_flushNext} != 2'b00) || ({writeback_arbitration_flushIt,{memaccess_arbitration_flushIt,execute_arbitration_flushIt}} != 3'b000));
  assign memaccess_arbitration_isFlushed = ((writeback_arbitration_flushNext != 1'b0) || ({writeback_arbitration_flushIt,memaccess_arbitration_flushIt} != 2'b00));
  assign writeback_arbitration_isFlushed = (1'b0 || (writeback_arbitration_flushIt != 1'b0));
  assign fetch_arbitration_isStuckByOthers = (fetch_arbitration_haltByOther || ((((1'b0 || decode_arbitration_isStuck) || execute_arbitration_isStuck) || memaccess_arbitration_isStuck) || writeback_arbitration_isStuck));
  assign fetch_arbitration_isStuck = (fetch_arbitration_haltItself || fetch_arbitration_isStuckByOthers);
  assign fetch_arbitration_isMoving = ((! fetch_arbitration_isStuck) && (! fetch_arbitration_removeIt));
  assign fetch_arbitration_isFiring = ((fetch_arbitration_isValid && (! fetch_arbitration_isStuck)) && (! fetch_arbitration_removeIt));
  assign decode_arbitration_isStuckByOthers = (decode_arbitration_haltByOther || (((1'b0 || execute_arbitration_isStuck) || memaccess_arbitration_isStuck) || writeback_arbitration_isStuck));
  assign decode_arbitration_isStuck = (decode_arbitration_haltItself || decode_arbitration_isStuckByOthers);
  assign decode_arbitration_isMoving = ((! decode_arbitration_isStuck) && (! decode_arbitration_removeIt));
  assign decode_arbitration_isFiring = ((decode_arbitration_isValid && (! decode_arbitration_isStuck)) && (! decode_arbitration_removeIt));
  assign execute_arbitration_isStuckByOthers = (execute_arbitration_haltByOther || ((1'b0 || memaccess_arbitration_isStuck) || writeback_arbitration_isStuck));
  assign execute_arbitration_isStuck = (execute_arbitration_haltItself || execute_arbitration_isStuckByOthers);
  assign execute_arbitration_isMoving = ((! execute_arbitration_isStuck) && (! execute_arbitration_removeIt));
  assign execute_arbitration_isFiring = ((execute_arbitration_isValid && (! execute_arbitration_isStuck)) && (! execute_arbitration_removeIt));
  assign memaccess_arbitration_isStuckByOthers = (memaccess_arbitration_haltByOther || (1'b0 || writeback_arbitration_isStuck));
  assign memaccess_arbitration_isStuck = (memaccess_arbitration_haltItself || memaccess_arbitration_isStuckByOthers);
  assign memaccess_arbitration_isMoving = ((! memaccess_arbitration_isStuck) && (! memaccess_arbitration_removeIt));
  assign memaccess_arbitration_isFiring = ((memaccess_arbitration_isValid && (! memaccess_arbitration_isStuck)) && (! memaccess_arbitration_removeIt));
  assign writeback_arbitration_isStuckByOthers = (writeback_arbitration_haltByOther || 1'b0);
  assign writeback_arbitration_isStuck = (writeback_arbitration_haltItself || writeback_arbitration_isStuckByOthers);
  assign writeback_arbitration_isMoving = ((! writeback_arbitration_isStuck) && (! writeback_arbitration_removeIt));
  assign writeback_arbitration_isFiring = ((writeback_arbitration_isValid && (! writeback_arbitration_isStuck)) && (! writeback_arbitration_removeIt));
  assign when_Pipeline_l163 = ((! fetch_arbitration_isStuck) && (! fetch_arbitration_removeIt));
  assign when_Pipeline_l166 = ((! decode_arbitration_isStuck) || decode_arbitration_removeIt);
  assign when_Pipeline_l163_1 = ((! decode_arbitration_isStuck) && (! decode_arbitration_removeIt));
  assign when_Pipeline_l166_1 = ((! execute_arbitration_isStuck) || execute_arbitration_removeIt);
  assign when_Pipeline_l163_2 = ((! execute_arbitration_isStuck) && (! execute_arbitration_removeIt));
  assign when_Pipeline_l166_2 = ((! memaccess_arbitration_isStuck) || memaccess_arbitration_removeIt);
  assign when_Pipeline_l163_3 = ((! memaccess_arbitration_isStuck) && (! memaccess_arbitration_removeIt));
  assign when_Pipeline_l166_3 = ((! writeback_arbitration_isStuck) || writeback_arbitration_removeIt);
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      pc_next <= 64'h0000000080000000;
      fetch_valid <= 1'b0;
      rsp_flush <= 1'b0;
      fetch_state <= IDLE;
      execute_ALUPlugin_branch_history <= 7'h0;
      _zz_when_DCachePlugin_l174 <= 1'b0;
      dcache_ar_valid <= 1'b0;
      dcache_ar_payload_id <= 4'b0000;
      dcache_ar_payload_len <= 8'h0;
      dcache_ar_payload_size <= 3'b000;
      dcache_ar_payload_burst <= 2'b00;
      dcache_ar_payload_addr <= 64'h0;
      dcache_aw_valid <= 1'b0;
      dcache_aw_payload_id <= 4'b0000;
      dcache_aw_payload_len <= 8'h0;
      dcache_aw_payload_size <= 3'b000;
      dcache_aw_payload_burst <= 2'b00;
      dcache_aw_payload_addr <= 64'h0;
      dcache_w_valid <= 1'b0;
      dcache_w_payload_data <= 64'h0;
      dcache_w_payload_strb <= 8'h0;
      dcache_w_payload_last <= 1'b0;
      decode_arbitration_isValid <= 1'b0;
      execute_arbitration_isValid <= 1'b0;
      memaccess_arbitration_isValid <= 1'b0;
      writeback_arbitration_isValid <= 1'b0;
    end else begin
      fetch_state <= fetch_state_next;
      if(when_FetchPlugin_l93) begin
        if(when_FetchPlugin_l94) begin
          rsp_flush <= 1'b1;
        end else begin
          if(when_FetchPlugin_l97) begin
            rsp_flush <= 1'b1;
          end else begin
            if(fetch_FetchPlugin_bpu_predict_taken) begin
              rsp_flush <= 1'b1;
            end
          end
        end
      end else begin
        if(ICachePlugin_icache_access_rsp_valid) begin
          rsp_flush <= 1'b0;
        end
      end
      if(when_FetchPlugin_l109) begin
        fetch_valid <= 1'b1;
      end else begin
        fetch_valid <= 1'b0;
      end
      if(when_FetchPlugin_l94) begin
        pc_next <= fetch_INT_PC;
      end else begin
        if(when_FetchPlugin_l97) begin
          pc_next <= _zz_pc_next;
        end else begin
          if(fetch_FetchPlugin_bpu_predict_taken) begin
            pc_next <= fetch_BPU_PC_NEXT;
          end else begin
            if(ICachePlugin_icache_access_cmd_fire_1) begin
              pc_next <= (pc_next + 64'h0000000000000004);
            end
          end
        end
      end
      if(execute_arbitration_isFiring) begin
        execute_ALUPlugin_branch_history <= {execute_ALUPlugin_branch_history[5 : 0],execute_ALUPlugin_branch_taken};
      end
      if(when_DCachePlugin_l118) begin
        dcache_ar_valid <= 1'b1;
      end else begin
        if(dcache_ar_fire) begin
          dcache_ar_valid <= 1'b0;
        end
      end
      dcache_ar_payload_id <= 4'b0001;
      dcache_ar_payload_len <= {4'd0, dCache_1_next_level_cmd_payload_len};
      dcache_ar_payload_size <= dCache_1_next_level_cmd_payload_size;
      dcache_ar_payload_burst <= 2'b01;
      dcache_ar_payload_addr <= dCache_1_next_level_cmd_payload_addr;
      if(when_DCachePlugin_l141) begin
        dcache_aw_valid <= 1'b1;
      end else begin
        if(dcache_aw_fire) begin
          dcache_aw_valid <= 1'b0;
        end
      end
      dcache_aw_payload_id <= 4'b0010;
      dcache_aw_payload_len <= {4'd0, dCache_1_next_level_cmd_payload_len};
      dcache_aw_payload_size <= dCache_1_next_level_cmd_payload_size;
      dcache_aw_payload_burst <= 2'b01;
      dcache_aw_payload_addr <= dCache_1_next_level_cmd_payload_addr;
      if(when_DCachePlugin_l159) begin
        dcache_w_valid <= 1'b1;
      end else begin
        if(dcache_w_fire) begin
          dcache_w_valid <= 1'b0;
        end
      end
      dcache_w_payload_data <= dCache_1_next_level_cmd_payload_wdata;
      dcache_w_payload_strb <= dCache_1_next_level_cmd_payload_wstrb;
      dcache_w_payload_last <= 1'b1;
      if(when_DCachePlugin_l174) begin
        if(when_DCachePlugin_l175) begin
          _zz_when_DCachePlugin_l174 <= 1'b0;
        end else begin
          if(when_DCachePlugin_l177) begin
            _zz_when_DCachePlugin_l174 <= 1'b1;
          end
        end
      end else begin
        if(when_DCachePlugin_l181) begin
          if(when_DCachePlugin_l182) begin
            _zz_when_DCachePlugin_l174 <= 1'b0;
          end
        end
      end
      if(when_Pipeline_l163) begin
        decode_arbitration_isValid <= fetch_arbitration_isValid;
      end else begin
        if(when_Pipeline_l166) begin
          decode_arbitration_isValid <= 1'b0;
        end
      end
      if(when_Pipeline_l163_1) begin
        execute_arbitration_isValid <= decode_arbitration_isValid;
      end else begin
        if(when_Pipeline_l166_1) begin
          execute_arbitration_isValid <= 1'b0;
        end
      end
      if(when_Pipeline_l163_2) begin
        memaccess_arbitration_isValid <= execute_arbitration_isValid;
      end else begin
        if(when_Pipeline_l166_2) begin
          memaccess_arbitration_isValid <= 1'b0;
        end
      end
      if(when_Pipeline_l163_3) begin
        writeback_arbitration_isValid <= memaccess_arbitration_isValid;
      end else begin
        if(when_Pipeline_l166_3) begin
          writeback_arbitration_isValid <= 1'b0;
        end
      end
    end
  end

  always @(posedge clk) begin
    if(when_Pipeline_l127) begin
      fetch_to_decode_PC <= fetch_PC;
    end
    if(when_Pipeline_l127_1) begin
      decode_to_execute_PC <= decode_PC;
    end
    if(when_Pipeline_l127_2) begin
      execute_to_memaccess_PC <= _zz_execute_to_memaccess_PC;
    end
    if(when_Pipeline_l127_3) begin
      memaccess_to_writeback_PC <= memaccess_PC;
    end
    if(when_Pipeline_l127_4) begin
      fetch_to_decode_PC_NEXT <= fetch_PC_NEXT;
    end
    if(when_Pipeline_l127_5) begin
      decode_to_execute_PC_NEXT <= decode_PC_NEXT;
    end
    if(when_Pipeline_l127_6) begin
      fetch_to_decode_INSTRUCTION <= fetch_INSTRUCTION;
    end
    if(when_Pipeline_l127_7) begin
      decode_to_execute_INSTRUCTION <= decode_INSTRUCTION;
    end
    if(when_Pipeline_l127_8) begin
      execute_to_memaccess_INSTRUCTION <= execute_INSTRUCTION;
    end
    if(when_Pipeline_l127_9) begin
      memaccess_to_writeback_INSTRUCTION <= memaccess_INSTRUCTION;
    end
    if(when_Pipeline_l127_10) begin
      fetch_to_decode_PREDICT_TAKEN <= fetch_PREDICT_TAKEN;
    end
    if(when_Pipeline_l127_11) begin
      decode_to_execute_PREDICT_TAKEN <= decode_PREDICT_TAKEN;
    end
    if(when_Pipeline_l127_12) begin
      decode_to_execute_IMM <= decode_IMM;
    end
    if(when_Pipeline_l127_13) begin
      decode_to_execute_RS1 <= decode_RS1;
    end
    if(when_Pipeline_l127_14) begin
      decode_to_execute_RS2 <= decode_RS2;
    end
    if(when_Pipeline_l127_15) begin
      decode_to_execute_RS1_ADDR <= decode_RS1_ADDR;
    end
    if(when_Pipeline_l127_16) begin
      decode_to_execute_RS2_ADDR <= decode_RS2_ADDR;
    end
    if(when_Pipeline_l127_17) begin
      decode_to_execute_ALU_CTRL <= decode_ALU_CTRL;
    end
    if(when_Pipeline_l127_18) begin
      decode_to_execute_ALU_WORD <= decode_ALU_WORD;
    end
    if(when_Pipeline_l127_19) begin
      decode_to_execute_SRC2_IS_IMM <= decode_SRC2_IS_IMM;
    end
    if(when_Pipeline_l127_20) begin
      decode_to_execute_MEM_CTRL <= decode_MEM_CTRL;
    end
    if(when_Pipeline_l127_21) begin
      execute_to_memaccess_MEM_CTRL <= execute_MEM_CTRL;
    end
    if(when_Pipeline_l127_22) begin
      decode_to_execute_RD_WEN <= decode_RD_WEN;
    end
    if(when_Pipeline_l127_23) begin
      execute_to_memaccess_RD_WEN <= execute_RD_WEN;
    end
    if(when_Pipeline_l127_24) begin
      memaccess_to_writeback_RD_WEN <= _zz_DecodePlugin_hazard_rs1_from_mem_3;
    end
    if(when_Pipeline_l127_25) begin
      decode_to_execute_RD_ADDR <= decode_RD_ADDR;
    end
    if(when_Pipeline_l127_26) begin
      execute_to_memaccess_RD_ADDR <= execute_RD_ADDR;
    end
    if(when_Pipeline_l127_27) begin
      memaccess_to_writeback_RD_ADDR <= _zz_DecodePlugin_hazard_rs1_from_mem_2;
    end
    if(when_Pipeline_l127_28) begin
      decode_to_execute_IS_LOAD <= decode_IS_LOAD;
    end
    if(when_Pipeline_l127_29) begin
      execute_to_memaccess_IS_LOAD <= execute_IS_LOAD;
    end
    if(when_Pipeline_l127_30) begin
      memaccess_to_writeback_IS_LOAD <= _zz_DecodePlugin_hazard_rs1_from_mem;
    end
    if(when_Pipeline_l127_31) begin
      decode_to_execute_IS_STORE <= decode_IS_STORE;
    end
    if(when_Pipeline_l127_32) begin
      execute_to_memaccess_IS_STORE <= execute_IS_STORE;
    end
    if(when_Pipeline_l127_33) begin
      decode_to_execute_CSR_CTRL <= decode_CSR_CTRL;
    end
    if(when_Pipeline_l127_34) begin
      decode_to_execute_CSR_ADDR <= _zz_decode_to_execute_CSR_ADDR;
    end
    if(when_Pipeline_l127_35) begin
      decode_to_execute_CSR_WEN <= decode_CSR_WEN;
    end
    if(when_Pipeline_l127_36) begin
      decode_to_execute_CSR_RDATA <= decode_CSR_RDATA;
    end
    if(when_Pipeline_l127_37) begin
      execute_to_memaccess_ALU_RESULT <= execute_ALU_RESULT;
    end
    if(when_Pipeline_l127_38) begin
      memaccess_to_writeback_ALU_RESULT <= _zz_execute_MEM_WDATA_1;
    end
    if(when_Pipeline_l127_39) begin
      execute_to_memaccess_MEM_WDATA <= execute_MEM_WDATA;
    end
    if(when_Pipeline_l127_40) begin
      memaccess_to_writeback_LSU_RDATA <= _zz_execute_MEM_WDATA;
    end
  end


endmodule

module SramBanks_1 (
  input               sram_0_ports_cmd_valid,
  input      [6:0]    sram_0_ports_cmd_payload_addr,
  input      [7:0]    sram_0_ports_cmd_payload_wen,
  input      [511:0]  sram_0_ports_cmd_payload_wdata,
  input      [63:0]   sram_0_ports_cmd_payload_wstrb,
  output              sram_0_ports_rsp_valid,
  output reg [511:0]  sram_0_ports_rsp_payload_data,
  input               sram_1_ports_cmd_valid,
  input      [6:0]    sram_1_ports_cmd_payload_addr,
  input      [7:0]    sram_1_ports_cmd_payload_wen,
  input      [511:0]  sram_1_ports_cmd_payload_wdata,
  input      [63:0]   sram_1_ports_cmd_payload_wstrb,
  output              sram_1_ports_rsp_valid,
  output reg [511:0]  sram_1_ports_rsp_payload_data,
  input               sram_2_ports_cmd_valid,
  input      [6:0]    sram_2_ports_cmd_payload_addr,
  input      [7:0]    sram_2_ports_cmd_payload_wen,
  input      [511:0]  sram_2_ports_cmd_payload_wdata,
  input      [63:0]   sram_2_ports_cmd_payload_wstrb,
  output              sram_2_ports_rsp_valid,
  output reg [511:0]  sram_2_ports_rsp_payload_data,
  input               sram_3_ports_cmd_valid,
  input      [6:0]    sram_3_ports_cmd_payload_addr,
  input      [7:0]    sram_3_ports_cmd_payload_wen,
  input      [511:0]  sram_3_ports_cmd_payload_wdata,
  input      [63:0]   sram_3_ports_cmd_payload_wstrb,
  output              sram_3_ports_rsp_valid,
  output reg [511:0]  sram_3_ports_rsp_payload_data,
  input               clk,
  input               reset
);

  wire       [63:0]   _zz_sram_0_banks_0_bank_port1;
  wire       [63:0]   _zz_sram_0_banks_1_bank_port1;
  wire       [63:0]   _zz_sram_0_banks_2_bank_port1;
  wire       [63:0]   _zz_sram_0_banks_3_bank_port1;
  wire       [63:0]   _zz_sram_0_banks_4_bank_port1;
  wire       [63:0]   _zz_sram_0_banks_5_bank_port1;
  wire       [63:0]   _zz_sram_0_banks_6_bank_port1;
  wire       [63:0]   _zz_sram_0_banks_7_bank_port1;
  wire       [63:0]   _zz_sram_1_banks_0_bank_port1;
  wire       [63:0]   _zz_sram_1_banks_1_bank_port1;
  wire       [63:0]   _zz_sram_1_banks_2_bank_port1;
  wire       [63:0]   _zz_sram_1_banks_3_bank_port1;
  wire       [63:0]   _zz_sram_1_banks_4_bank_port1;
  wire       [63:0]   _zz_sram_1_banks_5_bank_port1;
  wire       [63:0]   _zz_sram_1_banks_6_bank_port1;
  wire       [63:0]   _zz_sram_1_banks_7_bank_port1;
  wire       [63:0]   _zz_sram_2_banks_0_bank_port1;
  wire       [63:0]   _zz_sram_2_banks_1_bank_port1;
  wire       [63:0]   _zz_sram_2_banks_2_bank_port1;
  wire       [63:0]   _zz_sram_2_banks_3_bank_port1;
  wire       [63:0]   _zz_sram_2_banks_4_bank_port1;
  wire       [63:0]   _zz_sram_2_banks_5_bank_port1;
  wire       [63:0]   _zz_sram_2_banks_6_bank_port1;
  wire       [63:0]   _zz_sram_2_banks_7_bank_port1;
  wire       [63:0]   _zz_sram_3_banks_0_bank_port1;
  wire       [63:0]   _zz_sram_3_banks_1_bank_port1;
  wire       [63:0]   _zz_sram_3_banks_2_bank_port1;
  wire       [63:0]   _zz_sram_3_banks_3_bank_port1;
  wire       [63:0]   _zz_sram_3_banks_4_bank_port1;
  wire       [63:0]   _zz_sram_3_banks_5_bank_port1;
  wire       [63:0]   _zz_sram_3_banks_6_bank_port1;
  wire       [63:0]   _zz_sram_3_banks_7_bank_port1;
  wire       [63:0]   _zz_sram_0_banks_0_bank_port;
  wire       [7:0]    _zz_sram_0_banks_0_bank_port_1;
  wire                _zz_sram_0_banks_0_bank_port_2;
  wire       [63:0]   _zz_sram_0_banks_1_bank_port;
  wire       [7:0]    _zz_sram_0_banks_1_bank_port_1;
  wire                _zz_sram_0_banks_1_bank_port_2;
  wire       [63:0]   _zz_sram_0_banks_2_bank_port;
  wire       [7:0]    _zz_sram_0_banks_2_bank_port_1;
  wire                _zz_sram_0_banks_2_bank_port_2;
  wire       [63:0]   _zz_sram_0_banks_3_bank_port;
  wire       [7:0]    _zz_sram_0_banks_3_bank_port_1;
  wire                _zz_sram_0_banks_3_bank_port_2;
  wire       [63:0]   _zz_sram_0_banks_4_bank_port;
  wire       [7:0]    _zz_sram_0_banks_4_bank_port_1;
  wire                _zz_sram_0_banks_4_bank_port_2;
  wire       [63:0]   _zz_sram_0_banks_5_bank_port;
  wire       [7:0]    _zz_sram_0_banks_5_bank_port_1;
  wire                _zz_sram_0_banks_5_bank_port_2;
  wire       [63:0]   _zz_sram_0_banks_6_bank_port;
  wire       [7:0]    _zz_sram_0_banks_6_bank_port_1;
  wire                _zz_sram_0_banks_6_bank_port_2;
  wire       [63:0]   _zz_sram_0_banks_7_bank_port;
  wire       [7:0]    _zz_sram_0_banks_7_bank_port_1;
  wire                _zz_sram_0_banks_7_bank_port_2;
  wire       [63:0]   _zz_sram_1_banks_0_bank_port;
  wire       [7:0]    _zz_sram_1_banks_0_bank_port_1;
  wire                _zz_sram_1_banks_0_bank_port_2;
  wire       [63:0]   _zz_sram_1_banks_1_bank_port;
  wire       [7:0]    _zz_sram_1_banks_1_bank_port_1;
  wire                _zz_sram_1_banks_1_bank_port_2;
  wire       [63:0]   _zz_sram_1_banks_2_bank_port;
  wire       [7:0]    _zz_sram_1_banks_2_bank_port_1;
  wire                _zz_sram_1_banks_2_bank_port_2;
  wire       [63:0]   _zz_sram_1_banks_3_bank_port;
  wire       [7:0]    _zz_sram_1_banks_3_bank_port_1;
  wire                _zz_sram_1_banks_3_bank_port_2;
  wire       [63:0]   _zz_sram_1_banks_4_bank_port;
  wire       [7:0]    _zz_sram_1_banks_4_bank_port_1;
  wire                _zz_sram_1_banks_4_bank_port_2;
  wire       [63:0]   _zz_sram_1_banks_5_bank_port;
  wire       [7:0]    _zz_sram_1_banks_5_bank_port_1;
  wire                _zz_sram_1_banks_5_bank_port_2;
  wire       [63:0]   _zz_sram_1_banks_6_bank_port;
  wire       [7:0]    _zz_sram_1_banks_6_bank_port_1;
  wire                _zz_sram_1_banks_6_bank_port_2;
  wire       [63:0]   _zz_sram_1_banks_7_bank_port;
  wire       [7:0]    _zz_sram_1_banks_7_bank_port_1;
  wire                _zz_sram_1_banks_7_bank_port_2;
  wire       [63:0]   _zz_sram_2_banks_0_bank_port;
  wire       [7:0]    _zz_sram_2_banks_0_bank_port_1;
  wire                _zz_sram_2_banks_0_bank_port_2;
  wire       [63:0]   _zz_sram_2_banks_1_bank_port;
  wire       [7:0]    _zz_sram_2_banks_1_bank_port_1;
  wire                _zz_sram_2_banks_1_bank_port_2;
  wire       [63:0]   _zz_sram_2_banks_2_bank_port;
  wire       [7:0]    _zz_sram_2_banks_2_bank_port_1;
  wire                _zz_sram_2_banks_2_bank_port_2;
  wire       [63:0]   _zz_sram_2_banks_3_bank_port;
  wire       [7:0]    _zz_sram_2_banks_3_bank_port_1;
  wire                _zz_sram_2_banks_3_bank_port_2;
  wire       [63:0]   _zz_sram_2_banks_4_bank_port;
  wire       [7:0]    _zz_sram_2_banks_4_bank_port_1;
  wire                _zz_sram_2_banks_4_bank_port_2;
  wire       [63:0]   _zz_sram_2_banks_5_bank_port;
  wire       [7:0]    _zz_sram_2_banks_5_bank_port_1;
  wire                _zz_sram_2_banks_5_bank_port_2;
  wire       [63:0]   _zz_sram_2_banks_6_bank_port;
  wire       [7:0]    _zz_sram_2_banks_6_bank_port_1;
  wire                _zz_sram_2_banks_6_bank_port_2;
  wire       [63:0]   _zz_sram_2_banks_7_bank_port;
  wire       [7:0]    _zz_sram_2_banks_7_bank_port_1;
  wire                _zz_sram_2_banks_7_bank_port_2;
  wire       [63:0]   _zz_sram_3_banks_0_bank_port;
  wire       [7:0]    _zz_sram_3_banks_0_bank_port_1;
  wire                _zz_sram_3_banks_0_bank_port_2;
  wire       [63:0]   _zz_sram_3_banks_1_bank_port;
  wire       [7:0]    _zz_sram_3_banks_1_bank_port_1;
  wire                _zz_sram_3_banks_1_bank_port_2;
  wire       [63:0]   _zz_sram_3_banks_2_bank_port;
  wire       [7:0]    _zz_sram_3_banks_2_bank_port_1;
  wire                _zz_sram_3_banks_2_bank_port_2;
  wire       [63:0]   _zz_sram_3_banks_3_bank_port;
  wire       [7:0]    _zz_sram_3_banks_3_bank_port_1;
  wire                _zz_sram_3_banks_3_bank_port_2;
  wire       [63:0]   _zz_sram_3_banks_4_bank_port;
  wire       [7:0]    _zz_sram_3_banks_4_bank_port_1;
  wire                _zz_sram_3_banks_4_bank_port_2;
  wire       [63:0]   _zz_sram_3_banks_5_bank_port;
  wire       [7:0]    _zz_sram_3_banks_5_bank_port_1;
  wire                _zz_sram_3_banks_5_bank_port_2;
  wire       [63:0]   _zz_sram_3_banks_6_bank_port;
  wire       [7:0]    _zz_sram_3_banks_6_bank_port_1;
  wire                _zz_sram_3_banks_6_bank_port_2;
  wire       [63:0]   _zz_sram_3_banks_7_bank_port;
  wire       [7:0]    _zz_sram_3_banks_7_bank_port_1;
  wire                _zz_sram_3_banks_7_bank_port_2;
  reg                 _zz_sram_0_ports_rsp_valid;
  wire                when_SramBanks_l75;
  reg                 _zz_sram_1_ports_rsp_valid;
  wire                when_SramBanks_l75_1;
  reg                 _zz_sram_2_ports_rsp_valid;
  wire                when_SramBanks_l75_2;
  reg                 _zz_sram_3_ports_rsp_valid;
  wire                when_SramBanks_l75_3;
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_0_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_0_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_0_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_0_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_0_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_0_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_0_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_0_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_1_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_1_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_1_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_1_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_1_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_1_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_1_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_1_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_2_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_2_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_2_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_2_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_2_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_2_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_2_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_2_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_3_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_3_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_3_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_3_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_3_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_3_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_3_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_3_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_4_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_4_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_4_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_4_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_4_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_4_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_4_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_4_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_5_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_5_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_5_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_5_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_5_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_5_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_5_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_5_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_6_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_6_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_6_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_6_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_6_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_6_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_6_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_6_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_7_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_7_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_7_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_7_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_7_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_7_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_7_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_0_banks_7_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_0_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_0_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_0_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_0_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_0_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_0_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_0_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_0_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_1_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_1_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_1_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_1_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_1_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_1_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_1_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_1_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_2_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_2_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_2_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_2_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_2_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_2_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_2_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_2_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_3_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_3_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_3_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_3_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_3_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_3_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_3_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_3_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_4_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_4_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_4_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_4_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_4_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_4_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_4_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_4_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_5_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_5_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_5_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_5_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_5_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_5_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_5_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_5_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_6_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_6_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_6_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_6_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_6_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_6_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_6_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_6_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_7_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_7_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_7_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_7_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_7_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_7_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_7_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_1_banks_7_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_0_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_0_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_0_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_0_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_0_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_0_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_0_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_0_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_1_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_1_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_1_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_1_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_1_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_1_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_1_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_1_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_2_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_2_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_2_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_2_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_2_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_2_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_2_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_2_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_3_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_3_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_3_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_3_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_3_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_3_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_3_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_3_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_4_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_4_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_4_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_4_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_4_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_4_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_4_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_4_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_5_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_5_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_5_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_5_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_5_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_5_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_5_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_5_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_6_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_6_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_6_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_6_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_6_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_6_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_6_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_6_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_7_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_7_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_7_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_7_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_7_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_7_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_7_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_2_banks_7_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_0_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_0_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_0_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_0_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_0_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_0_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_0_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_0_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_1_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_1_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_1_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_1_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_1_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_1_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_1_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_1_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_2_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_2_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_2_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_2_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_2_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_2_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_2_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_2_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_3_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_3_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_3_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_3_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_3_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_3_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_3_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_3_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_4_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_4_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_4_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_4_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_4_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_4_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_4_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_4_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_5_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_5_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_5_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_5_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_5_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_5_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_5_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_5_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_6_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_6_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_6_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_6_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_6_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_6_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_6_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_6_bank_symbol7 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_7_bank_symbol0 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_7_bank_symbol1 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_7_bank_symbol2 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_7_bank_symbol3 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_7_bank_symbol4 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_7_bank_symbol5 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_7_bank_symbol6 [0:127];
  (* ram_style = "distributed" *) reg [7:0] sram_3_banks_7_bank_symbol7 [0:127];

  assign _zz_sram_0_banks_0_bank_port = sram_0_ports_cmd_payload_wdata[63 : 0];
  assign _zz_sram_0_banks_0_bank_port_1 = sram_0_ports_cmd_payload_wstrb[7 : 0];
  assign _zz_sram_0_banks_0_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[0]);
  assign _zz_sram_0_banks_1_bank_port = sram_0_ports_cmd_payload_wdata[127 : 64];
  assign _zz_sram_0_banks_1_bank_port_1 = sram_0_ports_cmd_payload_wstrb[15 : 8];
  assign _zz_sram_0_banks_1_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[1]);
  assign _zz_sram_0_banks_2_bank_port = sram_0_ports_cmd_payload_wdata[191 : 128];
  assign _zz_sram_0_banks_2_bank_port_1 = sram_0_ports_cmd_payload_wstrb[23 : 16];
  assign _zz_sram_0_banks_2_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[2]);
  assign _zz_sram_0_banks_3_bank_port = sram_0_ports_cmd_payload_wdata[255 : 192];
  assign _zz_sram_0_banks_3_bank_port_1 = sram_0_ports_cmd_payload_wstrb[31 : 24];
  assign _zz_sram_0_banks_3_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[3]);
  assign _zz_sram_0_banks_4_bank_port = sram_0_ports_cmd_payload_wdata[319 : 256];
  assign _zz_sram_0_banks_4_bank_port_1 = sram_0_ports_cmd_payload_wstrb[39 : 32];
  assign _zz_sram_0_banks_4_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[4]);
  assign _zz_sram_0_banks_5_bank_port = sram_0_ports_cmd_payload_wdata[383 : 320];
  assign _zz_sram_0_banks_5_bank_port_1 = sram_0_ports_cmd_payload_wstrb[47 : 40];
  assign _zz_sram_0_banks_5_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[5]);
  assign _zz_sram_0_banks_6_bank_port = sram_0_ports_cmd_payload_wdata[447 : 384];
  assign _zz_sram_0_banks_6_bank_port_1 = sram_0_ports_cmd_payload_wstrb[55 : 48];
  assign _zz_sram_0_banks_6_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[6]);
  assign _zz_sram_0_banks_7_bank_port = sram_0_ports_cmd_payload_wdata[511 : 448];
  assign _zz_sram_0_banks_7_bank_port_1 = sram_0_ports_cmd_payload_wstrb[63 : 56];
  assign _zz_sram_0_banks_7_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[7]);
  assign _zz_sram_1_banks_0_bank_port = sram_1_ports_cmd_payload_wdata[63 : 0];
  assign _zz_sram_1_banks_0_bank_port_1 = sram_1_ports_cmd_payload_wstrb[7 : 0];
  assign _zz_sram_1_banks_0_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[0]);
  assign _zz_sram_1_banks_1_bank_port = sram_1_ports_cmd_payload_wdata[127 : 64];
  assign _zz_sram_1_banks_1_bank_port_1 = sram_1_ports_cmd_payload_wstrb[15 : 8];
  assign _zz_sram_1_banks_1_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[1]);
  assign _zz_sram_1_banks_2_bank_port = sram_1_ports_cmd_payload_wdata[191 : 128];
  assign _zz_sram_1_banks_2_bank_port_1 = sram_1_ports_cmd_payload_wstrb[23 : 16];
  assign _zz_sram_1_banks_2_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[2]);
  assign _zz_sram_1_banks_3_bank_port = sram_1_ports_cmd_payload_wdata[255 : 192];
  assign _zz_sram_1_banks_3_bank_port_1 = sram_1_ports_cmd_payload_wstrb[31 : 24];
  assign _zz_sram_1_banks_3_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[3]);
  assign _zz_sram_1_banks_4_bank_port = sram_1_ports_cmd_payload_wdata[319 : 256];
  assign _zz_sram_1_banks_4_bank_port_1 = sram_1_ports_cmd_payload_wstrb[39 : 32];
  assign _zz_sram_1_banks_4_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[4]);
  assign _zz_sram_1_banks_5_bank_port = sram_1_ports_cmd_payload_wdata[383 : 320];
  assign _zz_sram_1_banks_5_bank_port_1 = sram_1_ports_cmd_payload_wstrb[47 : 40];
  assign _zz_sram_1_banks_5_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[5]);
  assign _zz_sram_1_banks_6_bank_port = sram_1_ports_cmd_payload_wdata[447 : 384];
  assign _zz_sram_1_banks_6_bank_port_1 = sram_1_ports_cmd_payload_wstrb[55 : 48];
  assign _zz_sram_1_banks_6_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[6]);
  assign _zz_sram_1_banks_7_bank_port = sram_1_ports_cmd_payload_wdata[511 : 448];
  assign _zz_sram_1_banks_7_bank_port_1 = sram_1_ports_cmd_payload_wstrb[63 : 56];
  assign _zz_sram_1_banks_7_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[7]);
  assign _zz_sram_2_banks_0_bank_port = sram_2_ports_cmd_payload_wdata[63 : 0];
  assign _zz_sram_2_banks_0_bank_port_1 = sram_2_ports_cmd_payload_wstrb[7 : 0];
  assign _zz_sram_2_banks_0_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[0]);
  assign _zz_sram_2_banks_1_bank_port = sram_2_ports_cmd_payload_wdata[127 : 64];
  assign _zz_sram_2_banks_1_bank_port_1 = sram_2_ports_cmd_payload_wstrb[15 : 8];
  assign _zz_sram_2_banks_1_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[1]);
  assign _zz_sram_2_banks_2_bank_port = sram_2_ports_cmd_payload_wdata[191 : 128];
  assign _zz_sram_2_banks_2_bank_port_1 = sram_2_ports_cmd_payload_wstrb[23 : 16];
  assign _zz_sram_2_banks_2_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[2]);
  assign _zz_sram_2_banks_3_bank_port = sram_2_ports_cmd_payload_wdata[255 : 192];
  assign _zz_sram_2_banks_3_bank_port_1 = sram_2_ports_cmd_payload_wstrb[31 : 24];
  assign _zz_sram_2_banks_3_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[3]);
  assign _zz_sram_2_banks_4_bank_port = sram_2_ports_cmd_payload_wdata[319 : 256];
  assign _zz_sram_2_banks_4_bank_port_1 = sram_2_ports_cmd_payload_wstrb[39 : 32];
  assign _zz_sram_2_banks_4_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[4]);
  assign _zz_sram_2_banks_5_bank_port = sram_2_ports_cmd_payload_wdata[383 : 320];
  assign _zz_sram_2_banks_5_bank_port_1 = sram_2_ports_cmd_payload_wstrb[47 : 40];
  assign _zz_sram_2_banks_5_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[5]);
  assign _zz_sram_2_banks_6_bank_port = sram_2_ports_cmd_payload_wdata[447 : 384];
  assign _zz_sram_2_banks_6_bank_port_1 = sram_2_ports_cmd_payload_wstrb[55 : 48];
  assign _zz_sram_2_banks_6_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[6]);
  assign _zz_sram_2_banks_7_bank_port = sram_2_ports_cmd_payload_wdata[511 : 448];
  assign _zz_sram_2_banks_7_bank_port_1 = sram_2_ports_cmd_payload_wstrb[63 : 56];
  assign _zz_sram_2_banks_7_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[7]);
  assign _zz_sram_3_banks_0_bank_port = sram_3_ports_cmd_payload_wdata[63 : 0];
  assign _zz_sram_3_banks_0_bank_port_1 = sram_3_ports_cmd_payload_wstrb[7 : 0];
  assign _zz_sram_3_banks_0_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[0]);
  assign _zz_sram_3_banks_1_bank_port = sram_3_ports_cmd_payload_wdata[127 : 64];
  assign _zz_sram_3_banks_1_bank_port_1 = sram_3_ports_cmd_payload_wstrb[15 : 8];
  assign _zz_sram_3_banks_1_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[1]);
  assign _zz_sram_3_banks_2_bank_port = sram_3_ports_cmd_payload_wdata[191 : 128];
  assign _zz_sram_3_banks_2_bank_port_1 = sram_3_ports_cmd_payload_wstrb[23 : 16];
  assign _zz_sram_3_banks_2_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[2]);
  assign _zz_sram_3_banks_3_bank_port = sram_3_ports_cmd_payload_wdata[255 : 192];
  assign _zz_sram_3_banks_3_bank_port_1 = sram_3_ports_cmd_payload_wstrb[31 : 24];
  assign _zz_sram_3_banks_3_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[3]);
  assign _zz_sram_3_banks_4_bank_port = sram_3_ports_cmd_payload_wdata[319 : 256];
  assign _zz_sram_3_banks_4_bank_port_1 = sram_3_ports_cmd_payload_wstrb[39 : 32];
  assign _zz_sram_3_banks_4_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[4]);
  assign _zz_sram_3_banks_5_bank_port = sram_3_ports_cmd_payload_wdata[383 : 320];
  assign _zz_sram_3_banks_5_bank_port_1 = sram_3_ports_cmd_payload_wstrb[47 : 40];
  assign _zz_sram_3_banks_5_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[5]);
  assign _zz_sram_3_banks_6_bank_port = sram_3_ports_cmd_payload_wdata[447 : 384];
  assign _zz_sram_3_banks_6_bank_port_1 = sram_3_ports_cmd_payload_wstrb[55 : 48];
  assign _zz_sram_3_banks_6_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[6]);
  assign _zz_sram_3_banks_7_bank_port = sram_3_ports_cmd_payload_wdata[511 : 448];
  assign _zz_sram_3_banks_7_bank_port_1 = sram_3_ports_cmd_payload_wstrb[63 : 56];
  assign _zz_sram_3_banks_7_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[7]);
  always @(posedge clk) begin
    if(_zz_sram_0_banks_0_bank_port_1[0] && _zz_sram_0_banks_0_bank_port_2) begin
      sram_0_banks_0_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_0_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_0_bank_port_1[1] && _zz_sram_0_banks_0_bank_port_2) begin
      sram_0_banks_0_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_0_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_0_bank_port_1[2] && _zz_sram_0_banks_0_bank_port_2) begin
      sram_0_banks_0_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_0_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_0_bank_port_1[3] && _zz_sram_0_banks_0_bank_port_2) begin
      sram_0_banks_0_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_0_bank_port[31 : 24];
    end
    if(_zz_sram_0_banks_0_bank_port_1[4] && _zz_sram_0_banks_0_bank_port_2) begin
      sram_0_banks_0_bank_symbol4[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_0_bank_port[39 : 32];
    end
    if(_zz_sram_0_banks_0_bank_port_1[5] && _zz_sram_0_banks_0_bank_port_2) begin
      sram_0_banks_0_bank_symbol5[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_0_bank_port[47 : 40];
    end
    if(_zz_sram_0_banks_0_bank_port_1[6] && _zz_sram_0_banks_0_bank_port_2) begin
      sram_0_banks_0_bank_symbol6[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_0_bank_port[55 : 48];
    end
    if(_zz_sram_0_banks_0_bank_port_1[7] && _zz_sram_0_banks_0_bank_port_2) begin
      sram_0_banks_0_bank_symbol7[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_0_bank_port[63 : 56];
    end
  end

  assign _zz_sram_0_banks_0_bank_port1[7 : 0] = sram_0_banks_0_bank_symbol0[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_0_bank_port1[15 : 8] = sram_0_banks_0_bank_symbol1[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_0_bank_port1[23 : 16] = sram_0_banks_0_bank_symbol2[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_0_bank_port1[31 : 24] = sram_0_banks_0_bank_symbol3[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_0_bank_port1[39 : 32] = sram_0_banks_0_bank_symbol4[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_0_bank_port1[47 : 40] = sram_0_banks_0_bank_symbol5[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_0_bank_port1[55 : 48] = sram_0_banks_0_bank_symbol6[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_0_bank_port1[63 : 56] = sram_0_banks_0_bank_symbol7[sram_0_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_0_banks_1_bank_port_1[0] && _zz_sram_0_banks_1_bank_port_2) begin
      sram_0_banks_1_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_1_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_1_bank_port_1[1] && _zz_sram_0_banks_1_bank_port_2) begin
      sram_0_banks_1_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_1_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_1_bank_port_1[2] && _zz_sram_0_banks_1_bank_port_2) begin
      sram_0_banks_1_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_1_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_1_bank_port_1[3] && _zz_sram_0_banks_1_bank_port_2) begin
      sram_0_banks_1_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_1_bank_port[31 : 24];
    end
    if(_zz_sram_0_banks_1_bank_port_1[4] && _zz_sram_0_banks_1_bank_port_2) begin
      sram_0_banks_1_bank_symbol4[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_1_bank_port[39 : 32];
    end
    if(_zz_sram_0_banks_1_bank_port_1[5] && _zz_sram_0_banks_1_bank_port_2) begin
      sram_0_banks_1_bank_symbol5[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_1_bank_port[47 : 40];
    end
    if(_zz_sram_0_banks_1_bank_port_1[6] && _zz_sram_0_banks_1_bank_port_2) begin
      sram_0_banks_1_bank_symbol6[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_1_bank_port[55 : 48];
    end
    if(_zz_sram_0_banks_1_bank_port_1[7] && _zz_sram_0_banks_1_bank_port_2) begin
      sram_0_banks_1_bank_symbol7[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_1_bank_port[63 : 56];
    end
  end

  assign _zz_sram_0_banks_1_bank_port1[7 : 0] = sram_0_banks_1_bank_symbol0[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_1_bank_port1[15 : 8] = sram_0_banks_1_bank_symbol1[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_1_bank_port1[23 : 16] = sram_0_banks_1_bank_symbol2[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_1_bank_port1[31 : 24] = sram_0_banks_1_bank_symbol3[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_1_bank_port1[39 : 32] = sram_0_banks_1_bank_symbol4[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_1_bank_port1[47 : 40] = sram_0_banks_1_bank_symbol5[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_1_bank_port1[55 : 48] = sram_0_banks_1_bank_symbol6[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_1_bank_port1[63 : 56] = sram_0_banks_1_bank_symbol7[sram_0_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_0_banks_2_bank_port_1[0] && _zz_sram_0_banks_2_bank_port_2) begin
      sram_0_banks_2_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_2_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_2_bank_port_1[1] && _zz_sram_0_banks_2_bank_port_2) begin
      sram_0_banks_2_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_2_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_2_bank_port_1[2] && _zz_sram_0_banks_2_bank_port_2) begin
      sram_0_banks_2_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_2_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_2_bank_port_1[3] && _zz_sram_0_banks_2_bank_port_2) begin
      sram_0_banks_2_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_2_bank_port[31 : 24];
    end
    if(_zz_sram_0_banks_2_bank_port_1[4] && _zz_sram_0_banks_2_bank_port_2) begin
      sram_0_banks_2_bank_symbol4[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_2_bank_port[39 : 32];
    end
    if(_zz_sram_0_banks_2_bank_port_1[5] && _zz_sram_0_banks_2_bank_port_2) begin
      sram_0_banks_2_bank_symbol5[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_2_bank_port[47 : 40];
    end
    if(_zz_sram_0_banks_2_bank_port_1[6] && _zz_sram_0_banks_2_bank_port_2) begin
      sram_0_banks_2_bank_symbol6[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_2_bank_port[55 : 48];
    end
    if(_zz_sram_0_banks_2_bank_port_1[7] && _zz_sram_0_banks_2_bank_port_2) begin
      sram_0_banks_2_bank_symbol7[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_2_bank_port[63 : 56];
    end
  end

  assign _zz_sram_0_banks_2_bank_port1[7 : 0] = sram_0_banks_2_bank_symbol0[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_2_bank_port1[15 : 8] = sram_0_banks_2_bank_symbol1[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_2_bank_port1[23 : 16] = sram_0_banks_2_bank_symbol2[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_2_bank_port1[31 : 24] = sram_0_banks_2_bank_symbol3[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_2_bank_port1[39 : 32] = sram_0_banks_2_bank_symbol4[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_2_bank_port1[47 : 40] = sram_0_banks_2_bank_symbol5[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_2_bank_port1[55 : 48] = sram_0_banks_2_bank_symbol6[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_2_bank_port1[63 : 56] = sram_0_banks_2_bank_symbol7[sram_0_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_0_banks_3_bank_port_1[0] && _zz_sram_0_banks_3_bank_port_2) begin
      sram_0_banks_3_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_3_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_3_bank_port_1[1] && _zz_sram_0_banks_3_bank_port_2) begin
      sram_0_banks_3_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_3_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_3_bank_port_1[2] && _zz_sram_0_banks_3_bank_port_2) begin
      sram_0_banks_3_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_3_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_3_bank_port_1[3] && _zz_sram_0_banks_3_bank_port_2) begin
      sram_0_banks_3_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_3_bank_port[31 : 24];
    end
    if(_zz_sram_0_banks_3_bank_port_1[4] && _zz_sram_0_banks_3_bank_port_2) begin
      sram_0_banks_3_bank_symbol4[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_3_bank_port[39 : 32];
    end
    if(_zz_sram_0_banks_3_bank_port_1[5] && _zz_sram_0_banks_3_bank_port_2) begin
      sram_0_banks_3_bank_symbol5[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_3_bank_port[47 : 40];
    end
    if(_zz_sram_0_banks_3_bank_port_1[6] && _zz_sram_0_banks_3_bank_port_2) begin
      sram_0_banks_3_bank_symbol6[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_3_bank_port[55 : 48];
    end
    if(_zz_sram_0_banks_3_bank_port_1[7] && _zz_sram_0_banks_3_bank_port_2) begin
      sram_0_banks_3_bank_symbol7[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_3_bank_port[63 : 56];
    end
  end

  assign _zz_sram_0_banks_3_bank_port1[7 : 0] = sram_0_banks_3_bank_symbol0[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_3_bank_port1[15 : 8] = sram_0_banks_3_bank_symbol1[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_3_bank_port1[23 : 16] = sram_0_banks_3_bank_symbol2[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_3_bank_port1[31 : 24] = sram_0_banks_3_bank_symbol3[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_3_bank_port1[39 : 32] = sram_0_banks_3_bank_symbol4[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_3_bank_port1[47 : 40] = sram_0_banks_3_bank_symbol5[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_3_bank_port1[55 : 48] = sram_0_banks_3_bank_symbol6[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_3_bank_port1[63 : 56] = sram_0_banks_3_bank_symbol7[sram_0_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_0_banks_4_bank_port_1[0] && _zz_sram_0_banks_4_bank_port_2) begin
      sram_0_banks_4_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_4_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_4_bank_port_1[1] && _zz_sram_0_banks_4_bank_port_2) begin
      sram_0_banks_4_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_4_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_4_bank_port_1[2] && _zz_sram_0_banks_4_bank_port_2) begin
      sram_0_banks_4_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_4_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_4_bank_port_1[3] && _zz_sram_0_banks_4_bank_port_2) begin
      sram_0_banks_4_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_4_bank_port[31 : 24];
    end
    if(_zz_sram_0_banks_4_bank_port_1[4] && _zz_sram_0_banks_4_bank_port_2) begin
      sram_0_banks_4_bank_symbol4[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_4_bank_port[39 : 32];
    end
    if(_zz_sram_0_banks_4_bank_port_1[5] && _zz_sram_0_banks_4_bank_port_2) begin
      sram_0_banks_4_bank_symbol5[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_4_bank_port[47 : 40];
    end
    if(_zz_sram_0_banks_4_bank_port_1[6] && _zz_sram_0_banks_4_bank_port_2) begin
      sram_0_banks_4_bank_symbol6[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_4_bank_port[55 : 48];
    end
    if(_zz_sram_0_banks_4_bank_port_1[7] && _zz_sram_0_banks_4_bank_port_2) begin
      sram_0_banks_4_bank_symbol7[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_4_bank_port[63 : 56];
    end
  end

  assign _zz_sram_0_banks_4_bank_port1[7 : 0] = sram_0_banks_4_bank_symbol0[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_4_bank_port1[15 : 8] = sram_0_banks_4_bank_symbol1[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_4_bank_port1[23 : 16] = sram_0_banks_4_bank_symbol2[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_4_bank_port1[31 : 24] = sram_0_banks_4_bank_symbol3[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_4_bank_port1[39 : 32] = sram_0_banks_4_bank_symbol4[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_4_bank_port1[47 : 40] = sram_0_banks_4_bank_symbol5[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_4_bank_port1[55 : 48] = sram_0_banks_4_bank_symbol6[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_4_bank_port1[63 : 56] = sram_0_banks_4_bank_symbol7[sram_0_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_0_banks_5_bank_port_1[0] && _zz_sram_0_banks_5_bank_port_2) begin
      sram_0_banks_5_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_5_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_5_bank_port_1[1] && _zz_sram_0_banks_5_bank_port_2) begin
      sram_0_banks_5_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_5_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_5_bank_port_1[2] && _zz_sram_0_banks_5_bank_port_2) begin
      sram_0_banks_5_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_5_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_5_bank_port_1[3] && _zz_sram_0_banks_5_bank_port_2) begin
      sram_0_banks_5_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_5_bank_port[31 : 24];
    end
    if(_zz_sram_0_banks_5_bank_port_1[4] && _zz_sram_0_banks_5_bank_port_2) begin
      sram_0_banks_5_bank_symbol4[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_5_bank_port[39 : 32];
    end
    if(_zz_sram_0_banks_5_bank_port_1[5] && _zz_sram_0_banks_5_bank_port_2) begin
      sram_0_banks_5_bank_symbol5[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_5_bank_port[47 : 40];
    end
    if(_zz_sram_0_banks_5_bank_port_1[6] && _zz_sram_0_banks_5_bank_port_2) begin
      sram_0_banks_5_bank_symbol6[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_5_bank_port[55 : 48];
    end
    if(_zz_sram_0_banks_5_bank_port_1[7] && _zz_sram_0_banks_5_bank_port_2) begin
      sram_0_banks_5_bank_symbol7[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_5_bank_port[63 : 56];
    end
  end

  assign _zz_sram_0_banks_5_bank_port1[7 : 0] = sram_0_banks_5_bank_symbol0[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_5_bank_port1[15 : 8] = sram_0_banks_5_bank_symbol1[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_5_bank_port1[23 : 16] = sram_0_banks_5_bank_symbol2[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_5_bank_port1[31 : 24] = sram_0_banks_5_bank_symbol3[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_5_bank_port1[39 : 32] = sram_0_banks_5_bank_symbol4[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_5_bank_port1[47 : 40] = sram_0_banks_5_bank_symbol5[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_5_bank_port1[55 : 48] = sram_0_banks_5_bank_symbol6[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_5_bank_port1[63 : 56] = sram_0_banks_5_bank_symbol7[sram_0_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_0_banks_6_bank_port_1[0] && _zz_sram_0_banks_6_bank_port_2) begin
      sram_0_banks_6_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_6_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_6_bank_port_1[1] && _zz_sram_0_banks_6_bank_port_2) begin
      sram_0_banks_6_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_6_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_6_bank_port_1[2] && _zz_sram_0_banks_6_bank_port_2) begin
      sram_0_banks_6_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_6_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_6_bank_port_1[3] && _zz_sram_0_banks_6_bank_port_2) begin
      sram_0_banks_6_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_6_bank_port[31 : 24];
    end
    if(_zz_sram_0_banks_6_bank_port_1[4] && _zz_sram_0_banks_6_bank_port_2) begin
      sram_0_banks_6_bank_symbol4[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_6_bank_port[39 : 32];
    end
    if(_zz_sram_0_banks_6_bank_port_1[5] && _zz_sram_0_banks_6_bank_port_2) begin
      sram_0_banks_6_bank_symbol5[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_6_bank_port[47 : 40];
    end
    if(_zz_sram_0_banks_6_bank_port_1[6] && _zz_sram_0_banks_6_bank_port_2) begin
      sram_0_banks_6_bank_symbol6[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_6_bank_port[55 : 48];
    end
    if(_zz_sram_0_banks_6_bank_port_1[7] && _zz_sram_0_banks_6_bank_port_2) begin
      sram_0_banks_6_bank_symbol7[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_6_bank_port[63 : 56];
    end
  end

  assign _zz_sram_0_banks_6_bank_port1[7 : 0] = sram_0_banks_6_bank_symbol0[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_6_bank_port1[15 : 8] = sram_0_banks_6_bank_symbol1[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_6_bank_port1[23 : 16] = sram_0_banks_6_bank_symbol2[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_6_bank_port1[31 : 24] = sram_0_banks_6_bank_symbol3[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_6_bank_port1[39 : 32] = sram_0_banks_6_bank_symbol4[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_6_bank_port1[47 : 40] = sram_0_banks_6_bank_symbol5[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_6_bank_port1[55 : 48] = sram_0_banks_6_bank_symbol6[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_6_bank_port1[63 : 56] = sram_0_banks_6_bank_symbol7[sram_0_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_0_banks_7_bank_port_1[0] && _zz_sram_0_banks_7_bank_port_2) begin
      sram_0_banks_7_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_7_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_7_bank_port_1[1] && _zz_sram_0_banks_7_bank_port_2) begin
      sram_0_banks_7_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_7_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_7_bank_port_1[2] && _zz_sram_0_banks_7_bank_port_2) begin
      sram_0_banks_7_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_7_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_7_bank_port_1[3] && _zz_sram_0_banks_7_bank_port_2) begin
      sram_0_banks_7_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_7_bank_port[31 : 24];
    end
    if(_zz_sram_0_banks_7_bank_port_1[4] && _zz_sram_0_banks_7_bank_port_2) begin
      sram_0_banks_7_bank_symbol4[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_7_bank_port[39 : 32];
    end
    if(_zz_sram_0_banks_7_bank_port_1[5] && _zz_sram_0_banks_7_bank_port_2) begin
      sram_0_banks_7_bank_symbol5[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_7_bank_port[47 : 40];
    end
    if(_zz_sram_0_banks_7_bank_port_1[6] && _zz_sram_0_banks_7_bank_port_2) begin
      sram_0_banks_7_bank_symbol6[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_7_bank_port[55 : 48];
    end
    if(_zz_sram_0_banks_7_bank_port_1[7] && _zz_sram_0_banks_7_bank_port_2) begin
      sram_0_banks_7_bank_symbol7[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_7_bank_port[63 : 56];
    end
  end

  assign _zz_sram_0_banks_7_bank_port1[7 : 0] = sram_0_banks_7_bank_symbol0[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_7_bank_port1[15 : 8] = sram_0_banks_7_bank_symbol1[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_7_bank_port1[23 : 16] = sram_0_banks_7_bank_symbol2[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_7_bank_port1[31 : 24] = sram_0_banks_7_bank_symbol3[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_7_bank_port1[39 : 32] = sram_0_banks_7_bank_symbol4[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_7_bank_port1[47 : 40] = sram_0_banks_7_bank_symbol5[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_7_bank_port1[55 : 48] = sram_0_banks_7_bank_symbol6[sram_0_ports_cmd_payload_addr];
  assign _zz_sram_0_banks_7_bank_port1[63 : 56] = sram_0_banks_7_bank_symbol7[sram_0_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_1_banks_0_bank_port_1[0] && _zz_sram_1_banks_0_bank_port_2) begin
      sram_1_banks_0_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_0_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_0_bank_port_1[1] && _zz_sram_1_banks_0_bank_port_2) begin
      sram_1_banks_0_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_0_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_0_bank_port_1[2] && _zz_sram_1_banks_0_bank_port_2) begin
      sram_1_banks_0_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_0_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_0_bank_port_1[3] && _zz_sram_1_banks_0_bank_port_2) begin
      sram_1_banks_0_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_0_bank_port[31 : 24];
    end
    if(_zz_sram_1_banks_0_bank_port_1[4] && _zz_sram_1_banks_0_bank_port_2) begin
      sram_1_banks_0_bank_symbol4[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_0_bank_port[39 : 32];
    end
    if(_zz_sram_1_banks_0_bank_port_1[5] && _zz_sram_1_banks_0_bank_port_2) begin
      sram_1_banks_0_bank_symbol5[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_0_bank_port[47 : 40];
    end
    if(_zz_sram_1_banks_0_bank_port_1[6] && _zz_sram_1_banks_0_bank_port_2) begin
      sram_1_banks_0_bank_symbol6[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_0_bank_port[55 : 48];
    end
    if(_zz_sram_1_banks_0_bank_port_1[7] && _zz_sram_1_banks_0_bank_port_2) begin
      sram_1_banks_0_bank_symbol7[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_0_bank_port[63 : 56];
    end
  end

  assign _zz_sram_1_banks_0_bank_port1[7 : 0] = sram_1_banks_0_bank_symbol0[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_0_bank_port1[15 : 8] = sram_1_banks_0_bank_symbol1[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_0_bank_port1[23 : 16] = sram_1_banks_0_bank_symbol2[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_0_bank_port1[31 : 24] = sram_1_banks_0_bank_symbol3[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_0_bank_port1[39 : 32] = sram_1_banks_0_bank_symbol4[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_0_bank_port1[47 : 40] = sram_1_banks_0_bank_symbol5[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_0_bank_port1[55 : 48] = sram_1_banks_0_bank_symbol6[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_0_bank_port1[63 : 56] = sram_1_banks_0_bank_symbol7[sram_1_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_1_banks_1_bank_port_1[0] && _zz_sram_1_banks_1_bank_port_2) begin
      sram_1_banks_1_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_1_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_1_bank_port_1[1] && _zz_sram_1_banks_1_bank_port_2) begin
      sram_1_banks_1_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_1_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_1_bank_port_1[2] && _zz_sram_1_banks_1_bank_port_2) begin
      sram_1_banks_1_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_1_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_1_bank_port_1[3] && _zz_sram_1_banks_1_bank_port_2) begin
      sram_1_banks_1_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_1_bank_port[31 : 24];
    end
    if(_zz_sram_1_banks_1_bank_port_1[4] && _zz_sram_1_banks_1_bank_port_2) begin
      sram_1_banks_1_bank_symbol4[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_1_bank_port[39 : 32];
    end
    if(_zz_sram_1_banks_1_bank_port_1[5] && _zz_sram_1_banks_1_bank_port_2) begin
      sram_1_banks_1_bank_symbol5[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_1_bank_port[47 : 40];
    end
    if(_zz_sram_1_banks_1_bank_port_1[6] && _zz_sram_1_banks_1_bank_port_2) begin
      sram_1_banks_1_bank_symbol6[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_1_bank_port[55 : 48];
    end
    if(_zz_sram_1_banks_1_bank_port_1[7] && _zz_sram_1_banks_1_bank_port_2) begin
      sram_1_banks_1_bank_symbol7[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_1_bank_port[63 : 56];
    end
  end

  assign _zz_sram_1_banks_1_bank_port1[7 : 0] = sram_1_banks_1_bank_symbol0[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_1_bank_port1[15 : 8] = sram_1_banks_1_bank_symbol1[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_1_bank_port1[23 : 16] = sram_1_banks_1_bank_symbol2[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_1_bank_port1[31 : 24] = sram_1_banks_1_bank_symbol3[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_1_bank_port1[39 : 32] = sram_1_banks_1_bank_symbol4[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_1_bank_port1[47 : 40] = sram_1_banks_1_bank_symbol5[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_1_bank_port1[55 : 48] = sram_1_banks_1_bank_symbol6[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_1_bank_port1[63 : 56] = sram_1_banks_1_bank_symbol7[sram_1_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_1_banks_2_bank_port_1[0] && _zz_sram_1_banks_2_bank_port_2) begin
      sram_1_banks_2_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_2_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_2_bank_port_1[1] && _zz_sram_1_banks_2_bank_port_2) begin
      sram_1_banks_2_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_2_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_2_bank_port_1[2] && _zz_sram_1_banks_2_bank_port_2) begin
      sram_1_banks_2_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_2_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_2_bank_port_1[3] && _zz_sram_1_banks_2_bank_port_2) begin
      sram_1_banks_2_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_2_bank_port[31 : 24];
    end
    if(_zz_sram_1_banks_2_bank_port_1[4] && _zz_sram_1_banks_2_bank_port_2) begin
      sram_1_banks_2_bank_symbol4[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_2_bank_port[39 : 32];
    end
    if(_zz_sram_1_banks_2_bank_port_1[5] && _zz_sram_1_banks_2_bank_port_2) begin
      sram_1_banks_2_bank_symbol5[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_2_bank_port[47 : 40];
    end
    if(_zz_sram_1_banks_2_bank_port_1[6] && _zz_sram_1_banks_2_bank_port_2) begin
      sram_1_banks_2_bank_symbol6[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_2_bank_port[55 : 48];
    end
    if(_zz_sram_1_banks_2_bank_port_1[7] && _zz_sram_1_banks_2_bank_port_2) begin
      sram_1_banks_2_bank_symbol7[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_2_bank_port[63 : 56];
    end
  end

  assign _zz_sram_1_banks_2_bank_port1[7 : 0] = sram_1_banks_2_bank_symbol0[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_2_bank_port1[15 : 8] = sram_1_banks_2_bank_symbol1[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_2_bank_port1[23 : 16] = sram_1_banks_2_bank_symbol2[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_2_bank_port1[31 : 24] = sram_1_banks_2_bank_symbol3[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_2_bank_port1[39 : 32] = sram_1_banks_2_bank_symbol4[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_2_bank_port1[47 : 40] = sram_1_banks_2_bank_symbol5[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_2_bank_port1[55 : 48] = sram_1_banks_2_bank_symbol6[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_2_bank_port1[63 : 56] = sram_1_banks_2_bank_symbol7[sram_1_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_1_banks_3_bank_port_1[0] && _zz_sram_1_banks_3_bank_port_2) begin
      sram_1_banks_3_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_3_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_3_bank_port_1[1] && _zz_sram_1_banks_3_bank_port_2) begin
      sram_1_banks_3_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_3_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_3_bank_port_1[2] && _zz_sram_1_banks_3_bank_port_2) begin
      sram_1_banks_3_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_3_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_3_bank_port_1[3] && _zz_sram_1_banks_3_bank_port_2) begin
      sram_1_banks_3_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_3_bank_port[31 : 24];
    end
    if(_zz_sram_1_banks_3_bank_port_1[4] && _zz_sram_1_banks_3_bank_port_2) begin
      sram_1_banks_3_bank_symbol4[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_3_bank_port[39 : 32];
    end
    if(_zz_sram_1_banks_3_bank_port_1[5] && _zz_sram_1_banks_3_bank_port_2) begin
      sram_1_banks_3_bank_symbol5[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_3_bank_port[47 : 40];
    end
    if(_zz_sram_1_banks_3_bank_port_1[6] && _zz_sram_1_banks_3_bank_port_2) begin
      sram_1_banks_3_bank_symbol6[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_3_bank_port[55 : 48];
    end
    if(_zz_sram_1_banks_3_bank_port_1[7] && _zz_sram_1_banks_3_bank_port_2) begin
      sram_1_banks_3_bank_symbol7[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_3_bank_port[63 : 56];
    end
  end

  assign _zz_sram_1_banks_3_bank_port1[7 : 0] = sram_1_banks_3_bank_symbol0[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_3_bank_port1[15 : 8] = sram_1_banks_3_bank_symbol1[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_3_bank_port1[23 : 16] = sram_1_banks_3_bank_symbol2[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_3_bank_port1[31 : 24] = sram_1_banks_3_bank_symbol3[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_3_bank_port1[39 : 32] = sram_1_banks_3_bank_symbol4[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_3_bank_port1[47 : 40] = sram_1_banks_3_bank_symbol5[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_3_bank_port1[55 : 48] = sram_1_banks_3_bank_symbol6[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_3_bank_port1[63 : 56] = sram_1_banks_3_bank_symbol7[sram_1_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_1_banks_4_bank_port_1[0] && _zz_sram_1_banks_4_bank_port_2) begin
      sram_1_banks_4_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_4_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_4_bank_port_1[1] && _zz_sram_1_banks_4_bank_port_2) begin
      sram_1_banks_4_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_4_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_4_bank_port_1[2] && _zz_sram_1_banks_4_bank_port_2) begin
      sram_1_banks_4_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_4_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_4_bank_port_1[3] && _zz_sram_1_banks_4_bank_port_2) begin
      sram_1_banks_4_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_4_bank_port[31 : 24];
    end
    if(_zz_sram_1_banks_4_bank_port_1[4] && _zz_sram_1_banks_4_bank_port_2) begin
      sram_1_banks_4_bank_symbol4[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_4_bank_port[39 : 32];
    end
    if(_zz_sram_1_banks_4_bank_port_1[5] && _zz_sram_1_banks_4_bank_port_2) begin
      sram_1_banks_4_bank_symbol5[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_4_bank_port[47 : 40];
    end
    if(_zz_sram_1_banks_4_bank_port_1[6] && _zz_sram_1_banks_4_bank_port_2) begin
      sram_1_banks_4_bank_symbol6[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_4_bank_port[55 : 48];
    end
    if(_zz_sram_1_banks_4_bank_port_1[7] && _zz_sram_1_banks_4_bank_port_2) begin
      sram_1_banks_4_bank_symbol7[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_4_bank_port[63 : 56];
    end
  end

  assign _zz_sram_1_banks_4_bank_port1[7 : 0] = sram_1_banks_4_bank_symbol0[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_4_bank_port1[15 : 8] = sram_1_banks_4_bank_symbol1[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_4_bank_port1[23 : 16] = sram_1_banks_4_bank_symbol2[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_4_bank_port1[31 : 24] = sram_1_banks_4_bank_symbol3[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_4_bank_port1[39 : 32] = sram_1_banks_4_bank_symbol4[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_4_bank_port1[47 : 40] = sram_1_banks_4_bank_symbol5[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_4_bank_port1[55 : 48] = sram_1_banks_4_bank_symbol6[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_4_bank_port1[63 : 56] = sram_1_banks_4_bank_symbol7[sram_1_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_1_banks_5_bank_port_1[0] && _zz_sram_1_banks_5_bank_port_2) begin
      sram_1_banks_5_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_5_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_5_bank_port_1[1] && _zz_sram_1_banks_5_bank_port_2) begin
      sram_1_banks_5_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_5_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_5_bank_port_1[2] && _zz_sram_1_banks_5_bank_port_2) begin
      sram_1_banks_5_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_5_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_5_bank_port_1[3] && _zz_sram_1_banks_5_bank_port_2) begin
      sram_1_banks_5_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_5_bank_port[31 : 24];
    end
    if(_zz_sram_1_banks_5_bank_port_1[4] && _zz_sram_1_banks_5_bank_port_2) begin
      sram_1_banks_5_bank_symbol4[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_5_bank_port[39 : 32];
    end
    if(_zz_sram_1_banks_5_bank_port_1[5] && _zz_sram_1_banks_5_bank_port_2) begin
      sram_1_banks_5_bank_symbol5[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_5_bank_port[47 : 40];
    end
    if(_zz_sram_1_banks_5_bank_port_1[6] && _zz_sram_1_banks_5_bank_port_2) begin
      sram_1_banks_5_bank_symbol6[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_5_bank_port[55 : 48];
    end
    if(_zz_sram_1_banks_5_bank_port_1[7] && _zz_sram_1_banks_5_bank_port_2) begin
      sram_1_banks_5_bank_symbol7[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_5_bank_port[63 : 56];
    end
  end

  assign _zz_sram_1_banks_5_bank_port1[7 : 0] = sram_1_banks_5_bank_symbol0[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_5_bank_port1[15 : 8] = sram_1_banks_5_bank_symbol1[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_5_bank_port1[23 : 16] = sram_1_banks_5_bank_symbol2[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_5_bank_port1[31 : 24] = sram_1_banks_5_bank_symbol3[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_5_bank_port1[39 : 32] = sram_1_banks_5_bank_symbol4[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_5_bank_port1[47 : 40] = sram_1_banks_5_bank_symbol5[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_5_bank_port1[55 : 48] = sram_1_banks_5_bank_symbol6[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_5_bank_port1[63 : 56] = sram_1_banks_5_bank_symbol7[sram_1_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_1_banks_6_bank_port_1[0] && _zz_sram_1_banks_6_bank_port_2) begin
      sram_1_banks_6_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_6_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_6_bank_port_1[1] && _zz_sram_1_banks_6_bank_port_2) begin
      sram_1_banks_6_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_6_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_6_bank_port_1[2] && _zz_sram_1_banks_6_bank_port_2) begin
      sram_1_banks_6_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_6_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_6_bank_port_1[3] && _zz_sram_1_banks_6_bank_port_2) begin
      sram_1_banks_6_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_6_bank_port[31 : 24];
    end
    if(_zz_sram_1_banks_6_bank_port_1[4] && _zz_sram_1_banks_6_bank_port_2) begin
      sram_1_banks_6_bank_symbol4[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_6_bank_port[39 : 32];
    end
    if(_zz_sram_1_banks_6_bank_port_1[5] && _zz_sram_1_banks_6_bank_port_2) begin
      sram_1_banks_6_bank_symbol5[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_6_bank_port[47 : 40];
    end
    if(_zz_sram_1_banks_6_bank_port_1[6] && _zz_sram_1_banks_6_bank_port_2) begin
      sram_1_banks_6_bank_symbol6[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_6_bank_port[55 : 48];
    end
    if(_zz_sram_1_banks_6_bank_port_1[7] && _zz_sram_1_banks_6_bank_port_2) begin
      sram_1_banks_6_bank_symbol7[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_6_bank_port[63 : 56];
    end
  end

  assign _zz_sram_1_banks_6_bank_port1[7 : 0] = sram_1_banks_6_bank_symbol0[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_6_bank_port1[15 : 8] = sram_1_banks_6_bank_symbol1[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_6_bank_port1[23 : 16] = sram_1_banks_6_bank_symbol2[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_6_bank_port1[31 : 24] = sram_1_banks_6_bank_symbol3[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_6_bank_port1[39 : 32] = sram_1_banks_6_bank_symbol4[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_6_bank_port1[47 : 40] = sram_1_banks_6_bank_symbol5[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_6_bank_port1[55 : 48] = sram_1_banks_6_bank_symbol6[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_6_bank_port1[63 : 56] = sram_1_banks_6_bank_symbol7[sram_1_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_1_banks_7_bank_port_1[0] && _zz_sram_1_banks_7_bank_port_2) begin
      sram_1_banks_7_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_7_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_7_bank_port_1[1] && _zz_sram_1_banks_7_bank_port_2) begin
      sram_1_banks_7_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_7_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_7_bank_port_1[2] && _zz_sram_1_banks_7_bank_port_2) begin
      sram_1_banks_7_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_7_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_7_bank_port_1[3] && _zz_sram_1_banks_7_bank_port_2) begin
      sram_1_banks_7_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_7_bank_port[31 : 24];
    end
    if(_zz_sram_1_banks_7_bank_port_1[4] && _zz_sram_1_banks_7_bank_port_2) begin
      sram_1_banks_7_bank_symbol4[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_7_bank_port[39 : 32];
    end
    if(_zz_sram_1_banks_7_bank_port_1[5] && _zz_sram_1_banks_7_bank_port_2) begin
      sram_1_banks_7_bank_symbol5[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_7_bank_port[47 : 40];
    end
    if(_zz_sram_1_banks_7_bank_port_1[6] && _zz_sram_1_banks_7_bank_port_2) begin
      sram_1_banks_7_bank_symbol6[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_7_bank_port[55 : 48];
    end
    if(_zz_sram_1_banks_7_bank_port_1[7] && _zz_sram_1_banks_7_bank_port_2) begin
      sram_1_banks_7_bank_symbol7[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_7_bank_port[63 : 56];
    end
  end

  assign _zz_sram_1_banks_7_bank_port1[7 : 0] = sram_1_banks_7_bank_symbol0[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_7_bank_port1[15 : 8] = sram_1_banks_7_bank_symbol1[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_7_bank_port1[23 : 16] = sram_1_banks_7_bank_symbol2[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_7_bank_port1[31 : 24] = sram_1_banks_7_bank_symbol3[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_7_bank_port1[39 : 32] = sram_1_banks_7_bank_symbol4[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_7_bank_port1[47 : 40] = sram_1_banks_7_bank_symbol5[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_7_bank_port1[55 : 48] = sram_1_banks_7_bank_symbol6[sram_1_ports_cmd_payload_addr];
  assign _zz_sram_1_banks_7_bank_port1[63 : 56] = sram_1_banks_7_bank_symbol7[sram_1_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_2_banks_0_bank_port_1[0] && _zz_sram_2_banks_0_bank_port_2) begin
      sram_2_banks_0_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_0_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_0_bank_port_1[1] && _zz_sram_2_banks_0_bank_port_2) begin
      sram_2_banks_0_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_0_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_0_bank_port_1[2] && _zz_sram_2_banks_0_bank_port_2) begin
      sram_2_banks_0_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_0_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_0_bank_port_1[3] && _zz_sram_2_banks_0_bank_port_2) begin
      sram_2_banks_0_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_0_bank_port[31 : 24];
    end
    if(_zz_sram_2_banks_0_bank_port_1[4] && _zz_sram_2_banks_0_bank_port_2) begin
      sram_2_banks_0_bank_symbol4[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_0_bank_port[39 : 32];
    end
    if(_zz_sram_2_banks_0_bank_port_1[5] && _zz_sram_2_banks_0_bank_port_2) begin
      sram_2_banks_0_bank_symbol5[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_0_bank_port[47 : 40];
    end
    if(_zz_sram_2_banks_0_bank_port_1[6] && _zz_sram_2_banks_0_bank_port_2) begin
      sram_2_banks_0_bank_symbol6[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_0_bank_port[55 : 48];
    end
    if(_zz_sram_2_banks_0_bank_port_1[7] && _zz_sram_2_banks_0_bank_port_2) begin
      sram_2_banks_0_bank_symbol7[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_0_bank_port[63 : 56];
    end
  end

  assign _zz_sram_2_banks_0_bank_port1[7 : 0] = sram_2_banks_0_bank_symbol0[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_0_bank_port1[15 : 8] = sram_2_banks_0_bank_symbol1[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_0_bank_port1[23 : 16] = sram_2_banks_0_bank_symbol2[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_0_bank_port1[31 : 24] = sram_2_banks_0_bank_symbol3[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_0_bank_port1[39 : 32] = sram_2_banks_0_bank_symbol4[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_0_bank_port1[47 : 40] = sram_2_banks_0_bank_symbol5[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_0_bank_port1[55 : 48] = sram_2_banks_0_bank_symbol6[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_0_bank_port1[63 : 56] = sram_2_banks_0_bank_symbol7[sram_2_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_2_banks_1_bank_port_1[0] && _zz_sram_2_banks_1_bank_port_2) begin
      sram_2_banks_1_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_1_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_1_bank_port_1[1] && _zz_sram_2_banks_1_bank_port_2) begin
      sram_2_banks_1_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_1_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_1_bank_port_1[2] && _zz_sram_2_banks_1_bank_port_2) begin
      sram_2_banks_1_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_1_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_1_bank_port_1[3] && _zz_sram_2_banks_1_bank_port_2) begin
      sram_2_banks_1_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_1_bank_port[31 : 24];
    end
    if(_zz_sram_2_banks_1_bank_port_1[4] && _zz_sram_2_banks_1_bank_port_2) begin
      sram_2_banks_1_bank_symbol4[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_1_bank_port[39 : 32];
    end
    if(_zz_sram_2_banks_1_bank_port_1[5] && _zz_sram_2_banks_1_bank_port_2) begin
      sram_2_banks_1_bank_symbol5[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_1_bank_port[47 : 40];
    end
    if(_zz_sram_2_banks_1_bank_port_1[6] && _zz_sram_2_banks_1_bank_port_2) begin
      sram_2_banks_1_bank_symbol6[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_1_bank_port[55 : 48];
    end
    if(_zz_sram_2_banks_1_bank_port_1[7] && _zz_sram_2_banks_1_bank_port_2) begin
      sram_2_banks_1_bank_symbol7[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_1_bank_port[63 : 56];
    end
  end

  assign _zz_sram_2_banks_1_bank_port1[7 : 0] = sram_2_banks_1_bank_symbol0[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_1_bank_port1[15 : 8] = sram_2_banks_1_bank_symbol1[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_1_bank_port1[23 : 16] = sram_2_banks_1_bank_symbol2[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_1_bank_port1[31 : 24] = sram_2_banks_1_bank_symbol3[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_1_bank_port1[39 : 32] = sram_2_banks_1_bank_symbol4[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_1_bank_port1[47 : 40] = sram_2_banks_1_bank_symbol5[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_1_bank_port1[55 : 48] = sram_2_banks_1_bank_symbol6[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_1_bank_port1[63 : 56] = sram_2_banks_1_bank_symbol7[sram_2_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_2_banks_2_bank_port_1[0] && _zz_sram_2_banks_2_bank_port_2) begin
      sram_2_banks_2_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_2_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_2_bank_port_1[1] && _zz_sram_2_banks_2_bank_port_2) begin
      sram_2_banks_2_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_2_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_2_bank_port_1[2] && _zz_sram_2_banks_2_bank_port_2) begin
      sram_2_banks_2_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_2_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_2_bank_port_1[3] && _zz_sram_2_banks_2_bank_port_2) begin
      sram_2_banks_2_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_2_bank_port[31 : 24];
    end
    if(_zz_sram_2_banks_2_bank_port_1[4] && _zz_sram_2_banks_2_bank_port_2) begin
      sram_2_banks_2_bank_symbol4[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_2_bank_port[39 : 32];
    end
    if(_zz_sram_2_banks_2_bank_port_1[5] && _zz_sram_2_banks_2_bank_port_2) begin
      sram_2_banks_2_bank_symbol5[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_2_bank_port[47 : 40];
    end
    if(_zz_sram_2_banks_2_bank_port_1[6] && _zz_sram_2_banks_2_bank_port_2) begin
      sram_2_banks_2_bank_symbol6[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_2_bank_port[55 : 48];
    end
    if(_zz_sram_2_banks_2_bank_port_1[7] && _zz_sram_2_banks_2_bank_port_2) begin
      sram_2_banks_2_bank_symbol7[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_2_bank_port[63 : 56];
    end
  end

  assign _zz_sram_2_banks_2_bank_port1[7 : 0] = sram_2_banks_2_bank_symbol0[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_2_bank_port1[15 : 8] = sram_2_banks_2_bank_symbol1[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_2_bank_port1[23 : 16] = sram_2_banks_2_bank_symbol2[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_2_bank_port1[31 : 24] = sram_2_banks_2_bank_symbol3[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_2_bank_port1[39 : 32] = sram_2_banks_2_bank_symbol4[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_2_bank_port1[47 : 40] = sram_2_banks_2_bank_symbol5[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_2_bank_port1[55 : 48] = sram_2_banks_2_bank_symbol6[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_2_bank_port1[63 : 56] = sram_2_banks_2_bank_symbol7[sram_2_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_2_banks_3_bank_port_1[0] && _zz_sram_2_banks_3_bank_port_2) begin
      sram_2_banks_3_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_3_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_3_bank_port_1[1] && _zz_sram_2_banks_3_bank_port_2) begin
      sram_2_banks_3_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_3_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_3_bank_port_1[2] && _zz_sram_2_banks_3_bank_port_2) begin
      sram_2_banks_3_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_3_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_3_bank_port_1[3] && _zz_sram_2_banks_3_bank_port_2) begin
      sram_2_banks_3_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_3_bank_port[31 : 24];
    end
    if(_zz_sram_2_banks_3_bank_port_1[4] && _zz_sram_2_banks_3_bank_port_2) begin
      sram_2_banks_3_bank_symbol4[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_3_bank_port[39 : 32];
    end
    if(_zz_sram_2_banks_3_bank_port_1[5] && _zz_sram_2_banks_3_bank_port_2) begin
      sram_2_banks_3_bank_symbol5[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_3_bank_port[47 : 40];
    end
    if(_zz_sram_2_banks_3_bank_port_1[6] && _zz_sram_2_banks_3_bank_port_2) begin
      sram_2_banks_3_bank_symbol6[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_3_bank_port[55 : 48];
    end
    if(_zz_sram_2_banks_3_bank_port_1[7] && _zz_sram_2_banks_3_bank_port_2) begin
      sram_2_banks_3_bank_symbol7[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_3_bank_port[63 : 56];
    end
  end

  assign _zz_sram_2_banks_3_bank_port1[7 : 0] = sram_2_banks_3_bank_symbol0[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_3_bank_port1[15 : 8] = sram_2_banks_3_bank_symbol1[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_3_bank_port1[23 : 16] = sram_2_banks_3_bank_symbol2[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_3_bank_port1[31 : 24] = sram_2_banks_3_bank_symbol3[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_3_bank_port1[39 : 32] = sram_2_banks_3_bank_symbol4[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_3_bank_port1[47 : 40] = sram_2_banks_3_bank_symbol5[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_3_bank_port1[55 : 48] = sram_2_banks_3_bank_symbol6[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_3_bank_port1[63 : 56] = sram_2_banks_3_bank_symbol7[sram_2_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_2_banks_4_bank_port_1[0] && _zz_sram_2_banks_4_bank_port_2) begin
      sram_2_banks_4_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_4_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_4_bank_port_1[1] && _zz_sram_2_banks_4_bank_port_2) begin
      sram_2_banks_4_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_4_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_4_bank_port_1[2] && _zz_sram_2_banks_4_bank_port_2) begin
      sram_2_banks_4_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_4_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_4_bank_port_1[3] && _zz_sram_2_banks_4_bank_port_2) begin
      sram_2_banks_4_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_4_bank_port[31 : 24];
    end
    if(_zz_sram_2_banks_4_bank_port_1[4] && _zz_sram_2_banks_4_bank_port_2) begin
      sram_2_banks_4_bank_symbol4[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_4_bank_port[39 : 32];
    end
    if(_zz_sram_2_banks_4_bank_port_1[5] && _zz_sram_2_banks_4_bank_port_2) begin
      sram_2_banks_4_bank_symbol5[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_4_bank_port[47 : 40];
    end
    if(_zz_sram_2_banks_4_bank_port_1[6] && _zz_sram_2_banks_4_bank_port_2) begin
      sram_2_banks_4_bank_symbol6[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_4_bank_port[55 : 48];
    end
    if(_zz_sram_2_banks_4_bank_port_1[7] && _zz_sram_2_banks_4_bank_port_2) begin
      sram_2_banks_4_bank_symbol7[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_4_bank_port[63 : 56];
    end
  end

  assign _zz_sram_2_banks_4_bank_port1[7 : 0] = sram_2_banks_4_bank_symbol0[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_4_bank_port1[15 : 8] = sram_2_banks_4_bank_symbol1[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_4_bank_port1[23 : 16] = sram_2_banks_4_bank_symbol2[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_4_bank_port1[31 : 24] = sram_2_banks_4_bank_symbol3[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_4_bank_port1[39 : 32] = sram_2_banks_4_bank_symbol4[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_4_bank_port1[47 : 40] = sram_2_banks_4_bank_symbol5[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_4_bank_port1[55 : 48] = sram_2_banks_4_bank_symbol6[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_4_bank_port1[63 : 56] = sram_2_banks_4_bank_symbol7[sram_2_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_2_banks_5_bank_port_1[0] && _zz_sram_2_banks_5_bank_port_2) begin
      sram_2_banks_5_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_5_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_5_bank_port_1[1] && _zz_sram_2_banks_5_bank_port_2) begin
      sram_2_banks_5_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_5_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_5_bank_port_1[2] && _zz_sram_2_banks_5_bank_port_2) begin
      sram_2_banks_5_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_5_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_5_bank_port_1[3] && _zz_sram_2_banks_5_bank_port_2) begin
      sram_2_banks_5_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_5_bank_port[31 : 24];
    end
    if(_zz_sram_2_banks_5_bank_port_1[4] && _zz_sram_2_banks_5_bank_port_2) begin
      sram_2_banks_5_bank_symbol4[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_5_bank_port[39 : 32];
    end
    if(_zz_sram_2_banks_5_bank_port_1[5] && _zz_sram_2_banks_5_bank_port_2) begin
      sram_2_banks_5_bank_symbol5[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_5_bank_port[47 : 40];
    end
    if(_zz_sram_2_banks_5_bank_port_1[6] && _zz_sram_2_banks_5_bank_port_2) begin
      sram_2_banks_5_bank_symbol6[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_5_bank_port[55 : 48];
    end
    if(_zz_sram_2_banks_5_bank_port_1[7] && _zz_sram_2_banks_5_bank_port_2) begin
      sram_2_banks_5_bank_symbol7[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_5_bank_port[63 : 56];
    end
  end

  assign _zz_sram_2_banks_5_bank_port1[7 : 0] = sram_2_banks_5_bank_symbol0[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_5_bank_port1[15 : 8] = sram_2_banks_5_bank_symbol1[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_5_bank_port1[23 : 16] = sram_2_banks_5_bank_symbol2[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_5_bank_port1[31 : 24] = sram_2_banks_5_bank_symbol3[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_5_bank_port1[39 : 32] = sram_2_banks_5_bank_symbol4[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_5_bank_port1[47 : 40] = sram_2_banks_5_bank_symbol5[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_5_bank_port1[55 : 48] = sram_2_banks_5_bank_symbol6[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_5_bank_port1[63 : 56] = sram_2_banks_5_bank_symbol7[sram_2_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_2_banks_6_bank_port_1[0] && _zz_sram_2_banks_6_bank_port_2) begin
      sram_2_banks_6_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_6_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_6_bank_port_1[1] && _zz_sram_2_banks_6_bank_port_2) begin
      sram_2_banks_6_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_6_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_6_bank_port_1[2] && _zz_sram_2_banks_6_bank_port_2) begin
      sram_2_banks_6_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_6_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_6_bank_port_1[3] && _zz_sram_2_banks_6_bank_port_2) begin
      sram_2_banks_6_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_6_bank_port[31 : 24];
    end
    if(_zz_sram_2_banks_6_bank_port_1[4] && _zz_sram_2_banks_6_bank_port_2) begin
      sram_2_banks_6_bank_symbol4[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_6_bank_port[39 : 32];
    end
    if(_zz_sram_2_banks_6_bank_port_1[5] && _zz_sram_2_banks_6_bank_port_2) begin
      sram_2_banks_6_bank_symbol5[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_6_bank_port[47 : 40];
    end
    if(_zz_sram_2_banks_6_bank_port_1[6] && _zz_sram_2_banks_6_bank_port_2) begin
      sram_2_banks_6_bank_symbol6[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_6_bank_port[55 : 48];
    end
    if(_zz_sram_2_banks_6_bank_port_1[7] && _zz_sram_2_banks_6_bank_port_2) begin
      sram_2_banks_6_bank_symbol7[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_6_bank_port[63 : 56];
    end
  end

  assign _zz_sram_2_banks_6_bank_port1[7 : 0] = sram_2_banks_6_bank_symbol0[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_6_bank_port1[15 : 8] = sram_2_banks_6_bank_symbol1[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_6_bank_port1[23 : 16] = sram_2_banks_6_bank_symbol2[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_6_bank_port1[31 : 24] = sram_2_banks_6_bank_symbol3[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_6_bank_port1[39 : 32] = sram_2_banks_6_bank_symbol4[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_6_bank_port1[47 : 40] = sram_2_banks_6_bank_symbol5[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_6_bank_port1[55 : 48] = sram_2_banks_6_bank_symbol6[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_6_bank_port1[63 : 56] = sram_2_banks_6_bank_symbol7[sram_2_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_2_banks_7_bank_port_1[0] && _zz_sram_2_banks_7_bank_port_2) begin
      sram_2_banks_7_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_7_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_7_bank_port_1[1] && _zz_sram_2_banks_7_bank_port_2) begin
      sram_2_banks_7_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_7_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_7_bank_port_1[2] && _zz_sram_2_banks_7_bank_port_2) begin
      sram_2_banks_7_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_7_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_7_bank_port_1[3] && _zz_sram_2_banks_7_bank_port_2) begin
      sram_2_banks_7_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_7_bank_port[31 : 24];
    end
    if(_zz_sram_2_banks_7_bank_port_1[4] && _zz_sram_2_banks_7_bank_port_2) begin
      sram_2_banks_7_bank_symbol4[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_7_bank_port[39 : 32];
    end
    if(_zz_sram_2_banks_7_bank_port_1[5] && _zz_sram_2_banks_7_bank_port_2) begin
      sram_2_banks_7_bank_symbol5[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_7_bank_port[47 : 40];
    end
    if(_zz_sram_2_banks_7_bank_port_1[6] && _zz_sram_2_banks_7_bank_port_2) begin
      sram_2_banks_7_bank_symbol6[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_7_bank_port[55 : 48];
    end
    if(_zz_sram_2_banks_7_bank_port_1[7] && _zz_sram_2_banks_7_bank_port_2) begin
      sram_2_banks_7_bank_symbol7[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_7_bank_port[63 : 56];
    end
  end

  assign _zz_sram_2_banks_7_bank_port1[7 : 0] = sram_2_banks_7_bank_symbol0[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_7_bank_port1[15 : 8] = sram_2_banks_7_bank_symbol1[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_7_bank_port1[23 : 16] = sram_2_banks_7_bank_symbol2[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_7_bank_port1[31 : 24] = sram_2_banks_7_bank_symbol3[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_7_bank_port1[39 : 32] = sram_2_banks_7_bank_symbol4[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_7_bank_port1[47 : 40] = sram_2_banks_7_bank_symbol5[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_7_bank_port1[55 : 48] = sram_2_banks_7_bank_symbol6[sram_2_ports_cmd_payload_addr];
  assign _zz_sram_2_banks_7_bank_port1[63 : 56] = sram_2_banks_7_bank_symbol7[sram_2_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_3_banks_0_bank_port_1[0] && _zz_sram_3_banks_0_bank_port_2) begin
      sram_3_banks_0_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_0_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_0_bank_port_1[1] && _zz_sram_3_banks_0_bank_port_2) begin
      sram_3_banks_0_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_0_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_0_bank_port_1[2] && _zz_sram_3_banks_0_bank_port_2) begin
      sram_3_banks_0_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_0_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_0_bank_port_1[3] && _zz_sram_3_banks_0_bank_port_2) begin
      sram_3_banks_0_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_0_bank_port[31 : 24];
    end
    if(_zz_sram_3_banks_0_bank_port_1[4] && _zz_sram_3_banks_0_bank_port_2) begin
      sram_3_banks_0_bank_symbol4[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_0_bank_port[39 : 32];
    end
    if(_zz_sram_3_banks_0_bank_port_1[5] && _zz_sram_3_banks_0_bank_port_2) begin
      sram_3_banks_0_bank_symbol5[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_0_bank_port[47 : 40];
    end
    if(_zz_sram_3_banks_0_bank_port_1[6] && _zz_sram_3_banks_0_bank_port_2) begin
      sram_3_banks_0_bank_symbol6[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_0_bank_port[55 : 48];
    end
    if(_zz_sram_3_banks_0_bank_port_1[7] && _zz_sram_3_banks_0_bank_port_2) begin
      sram_3_banks_0_bank_symbol7[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_0_bank_port[63 : 56];
    end
  end

  assign _zz_sram_3_banks_0_bank_port1[7 : 0] = sram_3_banks_0_bank_symbol0[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_0_bank_port1[15 : 8] = sram_3_banks_0_bank_symbol1[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_0_bank_port1[23 : 16] = sram_3_banks_0_bank_symbol2[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_0_bank_port1[31 : 24] = sram_3_banks_0_bank_symbol3[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_0_bank_port1[39 : 32] = sram_3_banks_0_bank_symbol4[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_0_bank_port1[47 : 40] = sram_3_banks_0_bank_symbol5[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_0_bank_port1[55 : 48] = sram_3_banks_0_bank_symbol6[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_0_bank_port1[63 : 56] = sram_3_banks_0_bank_symbol7[sram_3_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_3_banks_1_bank_port_1[0] && _zz_sram_3_banks_1_bank_port_2) begin
      sram_3_banks_1_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_1_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_1_bank_port_1[1] && _zz_sram_3_banks_1_bank_port_2) begin
      sram_3_banks_1_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_1_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_1_bank_port_1[2] && _zz_sram_3_banks_1_bank_port_2) begin
      sram_3_banks_1_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_1_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_1_bank_port_1[3] && _zz_sram_3_banks_1_bank_port_2) begin
      sram_3_banks_1_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_1_bank_port[31 : 24];
    end
    if(_zz_sram_3_banks_1_bank_port_1[4] && _zz_sram_3_banks_1_bank_port_2) begin
      sram_3_banks_1_bank_symbol4[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_1_bank_port[39 : 32];
    end
    if(_zz_sram_3_banks_1_bank_port_1[5] && _zz_sram_3_banks_1_bank_port_2) begin
      sram_3_banks_1_bank_symbol5[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_1_bank_port[47 : 40];
    end
    if(_zz_sram_3_banks_1_bank_port_1[6] && _zz_sram_3_banks_1_bank_port_2) begin
      sram_3_banks_1_bank_symbol6[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_1_bank_port[55 : 48];
    end
    if(_zz_sram_3_banks_1_bank_port_1[7] && _zz_sram_3_banks_1_bank_port_2) begin
      sram_3_banks_1_bank_symbol7[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_1_bank_port[63 : 56];
    end
  end

  assign _zz_sram_3_banks_1_bank_port1[7 : 0] = sram_3_banks_1_bank_symbol0[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_1_bank_port1[15 : 8] = sram_3_banks_1_bank_symbol1[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_1_bank_port1[23 : 16] = sram_3_banks_1_bank_symbol2[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_1_bank_port1[31 : 24] = sram_3_banks_1_bank_symbol3[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_1_bank_port1[39 : 32] = sram_3_banks_1_bank_symbol4[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_1_bank_port1[47 : 40] = sram_3_banks_1_bank_symbol5[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_1_bank_port1[55 : 48] = sram_3_banks_1_bank_symbol6[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_1_bank_port1[63 : 56] = sram_3_banks_1_bank_symbol7[sram_3_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_3_banks_2_bank_port_1[0] && _zz_sram_3_banks_2_bank_port_2) begin
      sram_3_banks_2_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_2_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_2_bank_port_1[1] && _zz_sram_3_banks_2_bank_port_2) begin
      sram_3_banks_2_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_2_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_2_bank_port_1[2] && _zz_sram_3_banks_2_bank_port_2) begin
      sram_3_banks_2_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_2_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_2_bank_port_1[3] && _zz_sram_3_banks_2_bank_port_2) begin
      sram_3_banks_2_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_2_bank_port[31 : 24];
    end
    if(_zz_sram_3_banks_2_bank_port_1[4] && _zz_sram_3_banks_2_bank_port_2) begin
      sram_3_banks_2_bank_symbol4[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_2_bank_port[39 : 32];
    end
    if(_zz_sram_3_banks_2_bank_port_1[5] && _zz_sram_3_banks_2_bank_port_2) begin
      sram_3_banks_2_bank_symbol5[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_2_bank_port[47 : 40];
    end
    if(_zz_sram_3_banks_2_bank_port_1[6] && _zz_sram_3_banks_2_bank_port_2) begin
      sram_3_banks_2_bank_symbol6[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_2_bank_port[55 : 48];
    end
    if(_zz_sram_3_banks_2_bank_port_1[7] && _zz_sram_3_banks_2_bank_port_2) begin
      sram_3_banks_2_bank_symbol7[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_2_bank_port[63 : 56];
    end
  end

  assign _zz_sram_3_banks_2_bank_port1[7 : 0] = sram_3_banks_2_bank_symbol0[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_2_bank_port1[15 : 8] = sram_3_banks_2_bank_symbol1[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_2_bank_port1[23 : 16] = sram_3_banks_2_bank_symbol2[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_2_bank_port1[31 : 24] = sram_3_banks_2_bank_symbol3[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_2_bank_port1[39 : 32] = sram_3_banks_2_bank_symbol4[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_2_bank_port1[47 : 40] = sram_3_banks_2_bank_symbol5[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_2_bank_port1[55 : 48] = sram_3_banks_2_bank_symbol6[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_2_bank_port1[63 : 56] = sram_3_banks_2_bank_symbol7[sram_3_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_3_banks_3_bank_port_1[0] && _zz_sram_3_banks_3_bank_port_2) begin
      sram_3_banks_3_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_3_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_3_bank_port_1[1] && _zz_sram_3_banks_3_bank_port_2) begin
      sram_3_banks_3_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_3_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_3_bank_port_1[2] && _zz_sram_3_banks_3_bank_port_2) begin
      sram_3_banks_3_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_3_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_3_bank_port_1[3] && _zz_sram_3_banks_3_bank_port_2) begin
      sram_3_banks_3_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_3_bank_port[31 : 24];
    end
    if(_zz_sram_3_banks_3_bank_port_1[4] && _zz_sram_3_banks_3_bank_port_2) begin
      sram_3_banks_3_bank_symbol4[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_3_bank_port[39 : 32];
    end
    if(_zz_sram_3_banks_3_bank_port_1[5] && _zz_sram_3_banks_3_bank_port_2) begin
      sram_3_banks_3_bank_symbol5[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_3_bank_port[47 : 40];
    end
    if(_zz_sram_3_banks_3_bank_port_1[6] && _zz_sram_3_banks_3_bank_port_2) begin
      sram_3_banks_3_bank_symbol6[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_3_bank_port[55 : 48];
    end
    if(_zz_sram_3_banks_3_bank_port_1[7] && _zz_sram_3_banks_3_bank_port_2) begin
      sram_3_banks_3_bank_symbol7[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_3_bank_port[63 : 56];
    end
  end

  assign _zz_sram_3_banks_3_bank_port1[7 : 0] = sram_3_banks_3_bank_symbol0[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_3_bank_port1[15 : 8] = sram_3_banks_3_bank_symbol1[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_3_bank_port1[23 : 16] = sram_3_banks_3_bank_symbol2[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_3_bank_port1[31 : 24] = sram_3_banks_3_bank_symbol3[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_3_bank_port1[39 : 32] = sram_3_banks_3_bank_symbol4[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_3_bank_port1[47 : 40] = sram_3_banks_3_bank_symbol5[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_3_bank_port1[55 : 48] = sram_3_banks_3_bank_symbol6[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_3_bank_port1[63 : 56] = sram_3_banks_3_bank_symbol7[sram_3_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_3_banks_4_bank_port_1[0] && _zz_sram_3_banks_4_bank_port_2) begin
      sram_3_banks_4_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_4_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_4_bank_port_1[1] && _zz_sram_3_banks_4_bank_port_2) begin
      sram_3_banks_4_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_4_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_4_bank_port_1[2] && _zz_sram_3_banks_4_bank_port_2) begin
      sram_3_banks_4_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_4_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_4_bank_port_1[3] && _zz_sram_3_banks_4_bank_port_2) begin
      sram_3_banks_4_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_4_bank_port[31 : 24];
    end
    if(_zz_sram_3_banks_4_bank_port_1[4] && _zz_sram_3_banks_4_bank_port_2) begin
      sram_3_banks_4_bank_symbol4[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_4_bank_port[39 : 32];
    end
    if(_zz_sram_3_banks_4_bank_port_1[5] && _zz_sram_3_banks_4_bank_port_2) begin
      sram_3_banks_4_bank_symbol5[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_4_bank_port[47 : 40];
    end
    if(_zz_sram_3_banks_4_bank_port_1[6] && _zz_sram_3_banks_4_bank_port_2) begin
      sram_3_banks_4_bank_symbol6[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_4_bank_port[55 : 48];
    end
    if(_zz_sram_3_banks_4_bank_port_1[7] && _zz_sram_3_banks_4_bank_port_2) begin
      sram_3_banks_4_bank_symbol7[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_4_bank_port[63 : 56];
    end
  end

  assign _zz_sram_3_banks_4_bank_port1[7 : 0] = sram_3_banks_4_bank_symbol0[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_4_bank_port1[15 : 8] = sram_3_banks_4_bank_symbol1[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_4_bank_port1[23 : 16] = sram_3_banks_4_bank_symbol2[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_4_bank_port1[31 : 24] = sram_3_banks_4_bank_symbol3[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_4_bank_port1[39 : 32] = sram_3_banks_4_bank_symbol4[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_4_bank_port1[47 : 40] = sram_3_banks_4_bank_symbol5[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_4_bank_port1[55 : 48] = sram_3_banks_4_bank_symbol6[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_4_bank_port1[63 : 56] = sram_3_banks_4_bank_symbol7[sram_3_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_3_banks_5_bank_port_1[0] && _zz_sram_3_banks_5_bank_port_2) begin
      sram_3_banks_5_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_5_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_5_bank_port_1[1] && _zz_sram_3_banks_5_bank_port_2) begin
      sram_3_banks_5_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_5_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_5_bank_port_1[2] && _zz_sram_3_banks_5_bank_port_2) begin
      sram_3_banks_5_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_5_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_5_bank_port_1[3] && _zz_sram_3_banks_5_bank_port_2) begin
      sram_3_banks_5_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_5_bank_port[31 : 24];
    end
    if(_zz_sram_3_banks_5_bank_port_1[4] && _zz_sram_3_banks_5_bank_port_2) begin
      sram_3_banks_5_bank_symbol4[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_5_bank_port[39 : 32];
    end
    if(_zz_sram_3_banks_5_bank_port_1[5] && _zz_sram_3_banks_5_bank_port_2) begin
      sram_3_banks_5_bank_symbol5[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_5_bank_port[47 : 40];
    end
    if(_zz_sram_3_banks_5_bank_port_1[6] && _zz_sram_3_banks_5_bank_port_2) begin
      sram_3_banks_5_bank_symbol6[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_5_bank_port[55 : 48];
    end
    if(_zz_sram_3_banks_5_bank_port_1[7] && _zz_sram_3_banks_5_bank_port_2) begin
      sram_3_banks_5_bank_symbol7[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_5_bank_port[63 : 56];
    end
  end

  assign _zz_sram_3_banks_5_bank_port1[7 : 0] = sram_3_banks_5_bank_symbol0[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_5_bank_port1[15 : 8] = sram_3_banks_5_bank_symbol1[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_5_bank_port1[23 : 16] = sram_3_banks_5_bank_symbol2[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_5_bank_port1[31 : 24] = sram_3_banks_5_bank_symbol3[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_5_bank_port1[39 : 32] = sram_3_banks_5_bank_symbol4[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_5_bank_port1[47 : 40] = sram_3_banks_5_bank_symbol5[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_5_bank_port1[55 : 48] = sram_3_banks_5_bank_symbol6[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_5_bank_port1[63 : 56] = sram_3_banks_5_bank_symbol7[sram_3_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_3_banks_6_bank_port_1[0] && _zz_sram_3_banks_6_bank_port_2) begin
      sram_3_banks_6_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_6_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_6_bank_port_1[1] && _zz_sram_3_banks_6_bank_port_2) begin
      sram_3_banks_6_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_6_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_6_bank_port_1[2] && _zz_sram_3_banks_6_bank_port_2) begin
      sram_3_banks_6_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_6_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_6_bank_port_1[3] && _zz_sram_3_banks_6_bank_port_2) begin
      sram_3_banks_6_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_6_bank_port[31 : 24];
    end
    if(_zz_sram_3_banks_6_bank_port_1[4] && _zz_sram_3_banks_6_bank_port_2) begin
      sram_3_banks_6_bank_symbol4[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_6_bank_port[39 : 32];
    end
    if(_zz_sram_3_banks_6_bank_port_1[5] && _zz_sram_3_banks_6_bank_port_2) begin
      sram_3_banks_6_bank_symbol5[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_6_bank_port[47 : 40];
    end
    if(_zz_sram_3_banks_6_bank_port_1[6] && _zz_sram_3_banks_6_bank_port_2) begin
      sram_3_banks_6_bank_symbol6[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_6_bank_port[55 : 48];
    end
    if(_zz_sram_3_banks_6_bank_port_1[7] && _zz_sram_3_banks_6_bank_port_2) begin
      sram_3_banks_6_bank_symbol7[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_6_bank_port[63 : 56];
    end
  end

  assign _zz_sram_3_banks_6_bank_port1[7 : 0] = sram_3_banks_6_bank_symbol0[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_6_bank_port1[15 : 8] = sram_3_banks_6_bank_symbol1[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_6_bank_port1[23 : 16] = sram_3_banks_6_bank_symbol2[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_6_bank_port1[31 : 24] = sram_3_banks_6_bank_symbol3[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_6_bank_port1[39 : 32] = sram_3_banks_6_bank_symbol4[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_6_bank_port1[47 : 40] = sram_3_banks_6_bank_symbol5[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_6_bank_port1[55 : 48] = sram_3_banks_6_bank_symbol6[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_6_bank_port1[63 : 56] = sram_3_banks_6_bank_symbol7[sram_3_ports_cmd_payload_addr];
  always @(posedge clk) begin
    if(_zz_sram_3_banks_7_bank_port_1[0] && _zz_sram_3_banks_7_bank_port_2) begin
      sram_3_banks_7_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_7_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_7_bank_port_1[1] && _zz_sram_3_banks_7_bank_port_2) begin
      sram_3_banks_7_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_7_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_7_bank_port_1[2] && _zz_sram_3_banks_7_bank_port_2) begin
      sram_3_banks_7_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_7_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_7_bank_port_1[3] && _zz_sram_3_banks_7_bank_port_2) begin
      sram_3_banks_7_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_7_bank_port[31 : 24];
    end
    if(_zz_sram_3_banks_7_bank_port_1[4] && _zz_sram_3_banks_7_bank_port_2) begin
      sram_3_banks_7_bank_symbol4[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_7_bank_port[39 : 32];
    end
    if(_zz_sram_3_banks_7_bank_port_1[5] && _zz_sram_3_banks_7_bank_port_2) begin
      sram_3_banks_7_bank_symbol5[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_7_bank_port[47 : 40];
    end
    if(_zz_sram_3_banks_7_bank_port_1[6] && _zz_sram_3_banks_7_bank_port_2) begin
      sram_3_banks_7_bank_symbol6[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_7_bank_port[55 : 48];
    end
    if(_zz_sram_3_banks_7_bank_port_1[7] && _zz_sram_3_banks_7_bank_port_2) begin
      sram_3_banks_7_bank_symbol7[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_7_bank_port[63 : 56];
    end
  end

  assign _zz_sram_3_banks_7_bank_port1[7 : 0] = sram_3_banks_7_bank_symbol0[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_7_bank_port1[15 : 8] = sram_3_banks_7_bank_symbol1[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_7_bank_port1[23 : 16] = sram_3_banks_7_bank_symbol2[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_7_bank_port1[31 : 24] = sram_3_banks_7_bank_symbol3[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_7_bank_port1[39 : 32] = sram_3_banks_7_bank_symbol4[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_7_bank_port1[47 : 40] = sram_3_banks_7_bank_symbol5[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_7_bank_port1[55 : 48] = sram_3_banks_7_bank_symbol6[sram_3_ports_cmd_payload_addr];
  assign _zz_sram_3_banks_7_bank_port1[63 : 56] = sram_3_banks_7_bank_symbol7[sram_3_ports_cmd_payload_addr];
  always @(*) begin
    sram_0_ports_rsp_payload_data[63 : 0] = _zz_sram_0_banks_0_bank_port1;
    sram_0_ports_rsp_payload_data[127 : 64] = _zz_sram_0_banks_1_bank_port1;
    sram_0_ports_rsp_payload_data[191 : 128] = _zz_sram_0_banks_2_bank_port1;
    sram_0_ports_rsp_payload_data[255 : 192] = _zz_sram_0_banks_3_bank_port1;
    sram_0_ports_rsp_payload_data[319 : 256] = _zz_sram_0_banks_4_bank_port1;
    sram_0_ports_rsp_payload_data[383 : 320] = _zz_sram_0_banks_5_bank_port1;
    sram_0_ports_rsp_payload_data[447 : 384] = _zz_sram_0_banks_6_bank_port1;
    sram_0_ports_rsp_payload_data[511 : 448] = _zz_sram_0_banks_7_bank_port1;
  end

  assign when_SramBanks_l75 = (sram_0_ports_cmd_valid && (sram_0_ports_cmd_payload_wen == 8'h0));
  always @(*) begin
    if(when_SramBanks_l75) begin
      _zz_sram_0_ports_rsp_valid = 1'b1;
    end else begin
      _zz_sram_0_ports_rsp_valid = 1'b0;
    end
  end

  assign sram_0_ports_rsp_valid = _zz_sram_0_ports_rsp_valid;
  always @(*) begin
    sram_1_ports_rsp_payload_data[63 : 0] = _zz_sram_1_banks_0_bank_port1;
    sram_1_ports_rsp_payload_data[127 : 64] = _zz_sram_1_banks_1_bank_port1;
    sram_1_ports_rsp_payload_data[191 : 128] = _zz_sram_1_banks_2_bank_port1;
    sram_1_ports_rsp_payload_data[255 : 192] = _zz_sram_1_banks_3_bank_port1;
    sram_1_ports_rsp_payload_data[319 : 256] = _zz_sram_1_banks_4_bank_port1;
    sram_1_ports_rsp_payload_data[383 : 320] = _zz_sram_1_banks_5_bank_port1;
    sram_1_ports_rsp_payload_data[447 : 384] = _zz_sram_1_banks_6_bank_port1;
    sram_1_ports_rsp_payload_data[511 : 448] = _zz_sram_1_banks_7_bank_port1;
  end

  assign when_SramBanks_l75_1 = (sram_1_ports_cmd_valid && (sram_1_ports_cmd_payload_wen == 8'h0));
  always @(*) begin
    if(when_SramBanks_l75_1) begin
      _zz_sram_1_ports_rsp_valid = 1'b1;
    end else begin
      _zz_sram_1_ports_rsp_valid = 1'b0;
    end
  end

  assign sram_1_ports_rsp_valid = _zz_sram_1_ports_rsp_valid;
  always @(*) begin
    sram_2_ports_rsp_payload_data[63 : 0] = _zz_sram_2_banks_0_bank_port1;
    sram_2_ports_rsp_payload_data[127 : 64] = _zz_sram_2_banks_1_bank_port1;
    sram_2_ports_rsp_payload_data[191 : 128] = _zz_sram_2_banks_2_bank_port1;
    sram_2_ports_rsp_payload_data[255 : 192] = _zz_sram_2_banks_3_bank_port1;
    sram_2_ports_rsp_payload_data[319 : 256] = _zz_sram_2_banks_4_bank_port1;
    sram_2_ports_rsp_payload_data[383 : 320] = _zz_sram_2_banks_5_bank_port1;
    sram_2_ports_rsp_payload_data[447 : 384] = _zz_sram_2_banks_6_bank_port1;
    sram_2_ports_rsp_payload_data[511 : 448] = _zz_sram_2_banks_7_bank_port1;
  end

  assign when_SramBanks_l75_2 = (sram_2_ports_cmd_valid && (sram_2_ports_cmd_payload_wen == 8'h0));
  always @(*) begin
    if(when_SramBanks_l75_2) begin
      _zz_sram_2_ports_rsp_valid = 1'b1;
    end else begin
      _zz_sram_2_ports_rsp_valid = 1'b0;
    end
  end

  assign sram_2_ports_rsp_valid = _zz_sram_2_ports_rsp_valid;
  always @(*) begin
    sram_3_ports_rsp_payload_data[63 : 0] = _zz_sram_3_banks_0_bank_port1;
    sram_3_ports_rsp_payload_data[127 : 64] = _zz_sram_3_banks_1_bank_port1;
    sram_3_ports_rsp_payload_data[191 : 128] = _zz_sram_3_banks_2_bank_port1;
    sram_3_ports_rsp_payload_data[255 : 192] = _zz_sram_3_banks_3_bank_port1;
    sram_3_ports_rsp_payload_data[319 : 256] = _zz_sram_3_banks_4_bank_port1;
    sram_3_ports_rsp_payload_data[383 : 320] = _zz_sram_3_banks_5_bank_port1;
    sram_3_ports_rsp_payload_data[447 : 384] = _zz_sram_3_banks_6_bank_port1;
    sram_3_ports_rsp_payload_data[511 : 448] = _zz_sram_3_banks_7_bank_port1;
  end

  assign when_SramBanks_l75_3 = (sram_3_ports_cmd_valid && (sram_3_ports_cmd_payload_wen == 8'h0));
  always @(*) begin
    if(when_SramBanks_l75_3) begin
      _zz_sram_3_ports_rsp_valid = 1'b1;
    end else begin
      _zz_sram_3_ports_rsp_valid = 1'b0;
    end
  end

  assign sram_3_ports_rsp_valid = _zz_sram_3_ports_rsp_valid;

endmodule

module DCache (
  output              stall,
  input               flush,
  input               cpu_cmd_valid,
  output              cpu_cmd_ready,
  input      [63:0]   cpu_cmd_payload_addr,
  input               cpu_cmd_payload_wen,
  input      [63:0]   cpu_cmd_payload_wdata,
  input      [7:0]    cpu_cmd_payload_wstrb,
  output              cpu_rsp_valid,
  output     [63:0]   cpu_rsp_payload_data,
  output reg          sram_0_ports_cmd_valid,
  output reg [6:0]    sram_0_ports_cmd_payload_addr,
  output reg [7:0]    sram_0_ports_cmd_payload_wen,
  output reg [511:0]  sram_0_ports_cmd_payload_wdata,
  output reg [63:0]   sram_0_ports_cmd_payload_wstrb,
  input               sram_0_ports_rsp_valid,
  input      [511:0]  sram_0_ports_rsp_payload_data,
  output reg          sram_1_ports_cmd_valid,
  output reg [6:0]    sram_1_ports_cmd_payload_addr,
  output reg [7:0]    sram_1_ports_cmd_payload_wen,
  output reg [511:0]  sram_1_ports_cmd_payload_wdata,
  output reg [63:0]   sram_1_ports_cmd_payload_wstrb,
  input               sram_1_ports_rsp_valid,
  input      [511:0]  sram_1_ports_rsp_payload_data,
  output reg          sram_2_ports_cmd_valid,
  output reg [6:0]    sram_2_ports_cmd_payload_addr,
  output reg [7:0]    sram_2_ports_cmd_payload_wen,
  output reg [511:0]  sram_2_ports_cmd_payload_wdata,
  output reg [63:0]   sram_2_ports_cmd_payload_wstrb,
  input               sram_2_ports_rsp_valid,
  input      [511:0]  sram_2_ports_rsp_payload_data,
  output reg          sram_3_ports_cmd_valid,
  output reg [6:0]    sram_3_ports_cmd_payload_addr,
  output reg [7:0]    sram_3_ports_cmd_payload_wen,
  output reg [511:0]  sram_3_ports_cmd_payload_wdata,
  output reg [63:0]   sram_3_ports_cmd_payload_wstrb,
  input               sram_3_ports_rsp_valid,
  input      [511:0]  sram_3_ports_rsp_payload_data,
  output              next_level_cmd_valid,
  input               next_level_cmd_ready,
  output     [63:0]   next_level_cmd_payload_addr,
  output     [3:0]    next_level_cmd_payload_len,
  output     [2:0]    next_level_cmd_payload_size,
  output              next_level_cmd_payload_wen,
  output     [63:0]   next_level_cmd_payload_wdata,
  output     [7:0]    next_level_cmd_payload_wstrb,
  input               next_level_rsp_valid,
  input      [63:0]   next_level_rsp_payload_data,
  input      [1:0]    next_level_rsp_payload_bresp,
  input               next_level_rsp_payload_rvalid,
  input               clk,
  input               reset
);

  wire       [6:0]    _zz_flush_cnt_valueNext;
  wire       [0:0]    _zz_flush_cnt_valueNext_1;
  wire       [2:0]    _zz_next_level_data_cnt_valueNext;
  wire       [0:0]    _zz_next_level_data_cnt_valueNext_1;
  wire       [6:0]    _zz_next_level_wstrb;
  wire       [7:0]    _zz__zz_cache_hit_gnt_0_3;
  wire       [7:0]    _zz__zz_cache_hit_gnt_0_3_1;
  wire       [3:0]    _zz__zz_cache_hit_gnt_0_3_2;
  wire       [7:0]    _zz__zz_cache_invld_gnt_0_3;
  wire       [7:0]    _zz__zz_cache_invld_gnt_0_3_1;
  wire       [3:0]    _zz__zz_cache_invld_gnt_0_3_2;
  wire       [7:0]    _zz__zz_cache_victim_gnt_0_3;
  wire       [7:0]    _zz__zz_cache_victim_gnt_0_3_1;
  wire       [3:0]    _zz__zz_cache_victim_gnt_0_3_2;
  reg                 _zz__zz_cache_hit_0;
  reg                 _zz__zz_cache_mru_0;
  reg        [50:0]   _zz_cache_tag_0;
  wire       [9:0]    _zz_sram_0_ports_cmd_payload_wdata;
  wire       [9:0]    _zz_sram_0_ports_cmd_payload_wstrb;
  wire       [9:0]    _zz_sram_0_ports_cmd_payload_wstrb_1;
  wire       [3:0]    _zz_sram_0_ports_cmd_payload_wen_1;
  wire       [9:0]    _zz_sram_0_ports_cmd_payload_wdata_1;
  wire       [9:0]    _zz_sram_0_ports_cmd_payload_wstrb_2;
  wire       [9:0]    _zz_sram_0_ports_cmd_payload_wstrb_3;
  reg                 _zz__zz_cache_hit_1;
  reg                 _zz__zz_cache_mru_1;
  reg        [50:0]   _zz_cache_tag_1;
  wire       [9:0]    _zz_sram_1_ports_cmd_payload_wdata;
  wire       [9:0]    _zz_sram_1_ports_cmd_payload_wstrb;
  wire       [9:0]    _zz_sram_1_ports_cmd_payload_wstrb_1;
  wire       [3:0]    _zz_sram_1_ports_cmd_payload_wen_1;
  wire       [9:0]    _zz_sram_1_ports_cmd_payload_wdata_1;
  wire       [9:0]    _zz_sram_1_ports_cmd_payload_wstrb_2;
  wire       [9:0]    _zz_sram_1_ports_cmd_payload_wstrb_3;
  reg                 _zz__zz_cache_hit_2;
  reg                 _zz__zz_cache_mru_2;
  reg        [50:0]   _zz_cache_tag_2;
  wire       [9:0]    _zz_sram_2_ports_cmd_payload_wdata;
  wire       [9:0]    _zz_sram_2_ports_cmd_payload_wstrb;
  wire       [9:0]    _zz_sram_2_ports_cmd_payload_wstrb_1;
  wire       [3:0]    _zz_sram_2_ports_cmd_payload_wen_1;
  wire       [9:0]    _zz_sram_2_ports_cmd_payload_wdata_1;
  wire       [9:0]    _zz_sram_2_ports_cmd_payload_wstrb_2;
  wire       [9:0]    _zz_sram_2_ports_cmd_payload_wstrb_3;
  reg                 _zz__zz_cache_hit_3;
  reg                 _zz__zz_cache_mru_3;
  reg        [50:0]   _zz_cache_tag_3;
  wire       [9:0]    _zz_sram_3_ports_cmd_payload_wdata;
  wire       [9:0]    _zz_sram_3_ports_cmd_payload_wstrb;
  wire       [9:0]    _zz_sram_3_ports_cmd_payload_wstrb_1;
  wire       [3:0]    _zz_sram_3_ports_cmd_payload_wen_1;
  wire       [9:0]    _zz_sram_3_ports_cmd_payload_wdata_1;
  wire       [9:0]    _zz_sram_3_ports_cmd_payload_wstrb_2;
  wire       [9:0]    _zz_sram_3_ports_cmd_payload_wstrb_3;
  reg        [511:0]  _zz__zz_cpu_rsp_payload_data;
  reg        [511:0]  _zz__zz_cpu_rsp_payload_data_1;
  reg        [63:0]   _zz_cpu_rsp_payload_data_2;
  reg        [63:0]   _zz_cpu_rsp_payload_data_3;
  reg                 _zz_cpu_rsp_valid;
  reg                 _zz_cpu_rsp_valid_1;
  wire                cpu_stall;
  reg                 ways_0_metas_0_vld;
  reg        [50:0]   ways_0_metas_0_tag;
  reg                 ways_0_metas_0_mru;
  reg                 ways_0_metas_1_vld;
  reg        [50:0]   ways_0_metas_1_tag;
  reg                 ways_0_metas_1_mru;
  reg                 ways_0_metas_2_vld;
  reg        [50:0]   ways_0_metas_2_tag;
  reg                 ways_0_metas_2_mru;
  reg                 ways_0_metas_3_vld;
  reg        [50:0]   ways_0_metas_3_tag;
  reg                 ways_0_metas_3_mru;
  reg                 ways_0_metas_4_vld;
  reg        [50:0]   ways_0_metas_4_tag;
  reg                 ways_0_metas_4_mru;
  reg                 ways_0_metas_5_vld;
  reg        [50:0]   ways_0_metas_5_tag;
  reg                 ways_0_metas_5_mru;
  reg                 ways_0_metas_6_vld;
  reg        [50:0]   ways_0_metas_6_tag;
  reg                 ways_0_metas_6_mru;
  reg                 ways_0_metas_7_vld;
  reg        [50:0]   ways_0_metas_7_tag;
  reg                 ways_0_metas_7_mru;
  reg                 ways_0_metas_8_vld;
  reg        [50:0]   ways_0_metas_8_tag;
  reg                 ways_0_metas_8_mru;
  reg                 ways_0_metas_9_vld;
  reg        [50:0]   ways_0_metas_9_tag;
  reg                 ways_0_metas_9_mru;
  reg                 ways_0_metas_10_vld;
  reg        [50:0]   ways_0_metas_10_tag;
  reg                 ways_0_metas_10_mru;
  reg                 ways_0_metas_11_vld;
  reg        [50:0]   ways_0_metas_11_tag;
  reg                 ways_0_metas_11_mru;
  reg                 ways_0_metas_12_vld;
  reg        [50:0]   ways_0_metas_12_tag;
  reg                 ways_0_metas_12_mru;
  reg                 ways_0_metas_13_vld;
  reg        [50:0]   ways_0_metas_13_tag;
  reg                 ways_0_metas_13_mru;
  reg                 ways_0_metas_14_vld;
  reg        [50:0]   ways_0_metas_14_tag;
  reg                 ways_0_metas_14_mru;
  reg                 ways_0_metas_15_vld;
  reg        [50:0]   ways_0_metas_15_tag;
  reg                 ways_0_metas_15_mru;
  reg                 ways_0_metas_16_vld;
  reg        [50:0]   ways_0_metas_16_tag;
  reg                 ways_0_metas_16_mru;
  reg                 ways_0_metas_17_vld;
  reg        [50:0]   ways_0_metas_17_tag;
  reg                 ways_0_metas_17_mru;
  reg                 ways_0_metas_18_vld;
  reg        [50:0]   ways_0_metas_18_tag;
  reg                 ways_0_metas_18_mru;
  reg                 ways_0_metas_19_vld;
  reg        [50:0]   ways_0_metas_19_tag;
  reg                 ways_0_metas_19_mru;
  reg                 ways_0_metas_20_vld;
  reg        [50:0]   ways_0_metas_20_tag;
  reg                 ways_0_metas_20_mru;
  reg                 ways_0_metas_21_vld;
  reg        [50:0]   ways_0_metas_21_tag;
  reg                 ways_0_metas_21_mru;
  reg                 ways_0_metas_22_vld;
  reg        [50:0]   ways_0_metas_22_tag;
  reg                 ways_0_metas_22_mru;
  reg                 ways_0_metas_23_vld;
  reg        [50:0]   ways_0_metas_23_tag;
  reg                 ways_0_metas_23_mru;
  reg                 ways_0_metas_24_vld;
  reg        [50:0]   ways_0_metas_24_tag;
  reg                 ways_0_metas_24_mru;
  reg                 ways_0_metas_25_vld;
  reg        [50:0]   ways_0_metas_25_tag;
  reg                 ways_0_metas_25_mru;
  reg                 ways_0_metas_26_vld;
  reg        [50:0]   ways_0_metas_26_tag;
  reg                 ways_0_metas_26_mru;
  reg                 ways_0_metas_27_vld;
  reg        [50:0]   ways_0_metas_27_tag;
  reg                 ways_0_metas_27_mru;
  reg                 ways_0_metas_28_vld;
  reg        [50:0]   ways_0_metas_28_tag;
  reg                 ways_0_metas_28_mru;
  reg                 ways_0_metas_29_vld;
  reg        [50:0]   ways_0_metas_29_tag;
  reg                 ways_0_metas_29_mru;
  reg                 ways_0_metas_30_vld;
  reg        [50:0]   ways_0_metas_30_tag;
  reg                 ways_0_metas_30_mru;
  reg                 ways_0_metas_31_vld;
  reg        [50:0]   ways_0_metas_31_tag;
  reg                 ways_0_metas_31_mru;
  reg                 ways_0_metas_32_vld;
  reg        [50:0]   ways_0_metas_32_tag;
  reg                 ways_0_metas_32_mru;
  reg                 ways_0_metas_33_vld;
  reg        [50:0]   ways_0_metas_33_tag;
  reg                 ways_0_metas_33_mru;
  reg                 ways_0_metas_34_vld;
  reg        [50:0]   ways_0_metas_34_tag;
  reg                 ways_0_metas_34_mru;
  reg                 ways_0_metas_35_vld;
  reg        [50:0]   ways_0_metas_35_tag;
  reg                 ways_0_metas_35_mru;
  reg                 ways_0_metas_36_vld;
  reg        [50:0]   ways_0_metas_36_tag;
  reg                 ways_0_metas_36_mru;
  reg                 ways_0_metas_37_vld;
  reg        [50:0]   ways_0_metas_37_tag;
  reg                 ways_0_metas_37_mru;
  reg                 ways_0_metas_38_vld;
  reg        [50:0]   ways_0_metas_38_tag;
  reg                 ways_0_metas_38_mru;
  reg                 ways_0_metas_39_vld;
  reg        [50:0]   ways_0_metas_39_tag;
  reg                 ways_0_metas_39_mru;
  reg                 ways_0_metas_40_vld;
  reg        [50:0]   ways_0_metas_40_tag;
  reg                 ways_0_metas_40_mru;
  reg                 ways_0_metas_41_vld;
  reg        [50:0]   ways_0_metas_41_tag;
  reg                 ways_0_metas_41_mru;
  reg                 ways_0_metas_42_vld;
  reg        [50:0]   ways_0_metas_42_tag;
  reg                 ways_0_metas_42_mru;
  reg                 ways_0_metas_43_vld;
  reg        [50:0]   ways_0_metas_43_tag;
  reg                 ways_0_metas_43_mru;
  reg                 ways_0_metas_44_vld;
  reg        [50:0]   ways_0_metas_44_tag;
  reg                 ways_0_metas_44_mru;
  reg                 ways_0_metas_45_vld;
  reg        [50:0]   ways_0_metas_45_tag;
  reg                 ways_0_metas_45_mru;
  reg                 ways_0_metas_46_vld;
  reg        [50:0]   ways_0_metas_46_tag;
  reg                 ways_0_metas_46_mru;
  reg                 ways_0_metas_47_vld;
  reg        [50:0]   ways_0_metas_47_tag;
  reg                 ways_0_metas_47_mru;
  reg                 ways_0_metas_48_vld;
  reg        [50:0]   ways_0_metas_48_tag;
  reg                 ways_0_metas_48_mru;
  reg                 ways_0_metas_49_vld;
  reg        [50:0]   ways_0_metas_49_tag;
  reg                 ways_0_metas_49_mru;
  reg                 ways_0_metas_50_vld;
  reg        [50:0]   ways_0_metas_50_tag;
  reg                 ways_0_metas_50_mru;
  reg                 ways_0_metas_51_vld;
  reg        [50:0]   ways_0_metas_51_tag;
  reg                 ways_0_metas_51_mru;
  reg                 ways_0_metas_52_vld;
  reg        [50:0]   ways_0_metas_52_tag;
  reg                 ways_0_metas_52_mru;
  reg                 ways_0_metas_53_vld;
  reg        [50:0]   ways_0_metas_53_tag;
  reg                 ways_0_metas_53_mru;
  reg                 ways_0_metas_54_vld;
  reg        [50:0]   ways_0_metas_54_tag;
  reg                 ways_0_metas_54_mru;
  reg                 ways_0_metas_55_vld;
  reg        [50:0]   ways_0_metas_55_tag;
  reg                 ways_0_metas_55_mru;
  reg                 ways_0_metas_56_vld;
  reg        [50:0]   ways_0_metas_56_tag;
  reg                 ways_0_metas_56_mru;
  reg                 ways_0_metas_57_vld;
  reg        [50:0]   ways_0_metas_57_tag;
  reg                 ways_0_metas_57_mru;
  reg                 ways_0_metas_58_vld;
  reg        [50:0]   ways_0_metas_58_tag;
  reg                 ways_0_metas_58_mru;
  reg                 ways_0_metas_59_vld;
  reg        [50:0]   ways_0_metas_59_tag;
  reg                 ways_0_metas_59_mru;
  reg                 ways_0_metas_60_vld;
  reg        [50:0]   ways_0_metas_60_tag;
  reg                 ways_0_metas_60_mru;
  reg                 ways_0_metas_61_vld;
  reg        [50:0]   ways_0_metas_61_tag;
  reg                 ways_0_metas_61_mru;
  reg                 ways_0_metas_62_vld;
  reg        [50:0]   ways_0_metas_62_tag;
  reg                 ways_0_metas_62_mru;
  reg                 ways_0_metas_63_vld;
  reg        [50:0]   ways_0_metas_63_tag;
  reg                 ways_0_metas_63_mru;
  reg                 ways_0_metas_64_vld;
  reg        [50:0]   ways_0_metas_64_tag;
  reg                 ways_0_metas_64_mru;
  reg                 ways_0_metas_65_vld;
  reg        [50:0]   ways_0_metas_65_tag;
  reg                 ways_0_metas_65_mru;
  reg                 ways_0_metas_66_vld;
  reg        [50:0]   ways_0_metas_66_tag;
  reg                 ways_0_metas_66_mru;
  reg                 ways_0_metas_67_vld;
  reg        [50:0]   ways_0_metas_67_tag;
  reg                 ways_0_metas_67_mru;
  reg                 ways_0_metas_68_vld;
  reg        [50:0]   ways_0_metas_68_tag;
  reg                 ways_0_metas_68_mru;
  reg                 ways_0_metas_69_vld;
  reg        [50:0]   ways_0_metas_69_tag;
  reg                 ways_0_metas_69_mru;
  reg                 ways_0_metas_70_vld;
  reg        [50:0]   ways_0_metas_70_tag;
  reg                 ways_0_metas_70_mru;
  reg                 ways_0_metas_71_vld;
  reg        [50:0]   ways_0_metas_71_tag;
  reg                 ways_0_metas_71_mru;
  reg                 ways_0_metas_72_vld;
  reg        [50:0]   ways_0_metas_72_tag;
  reg                 ways_0_metas_72_mru;
  reg                 ways_0_metas_73_vld;
  reg        [50:0]   ways_0_metas_73_tag;
  reg                 ways_0_metas_73_mru;
  reg                 ways_0_metas_74_vld;
  reg        [50:0]   ways_0_metas_74_tag;
  reg                 ways_0_metas_74_mru;
  reg                 ways_0_metas_75_vld;
  reg        [50:0]   ways_0_metas_75_tag;
  reg                 ways_0_metas_75_mru;
  reg                 ways_0_metas_76_vld;
  reg        [50:0]   ways_0_metas_76_tag;
  reg                 ways_0_metas_76_mru;
  reg                 ways_0_metas_77_vld;
  reg        [50:0]   ways_0_metas_77_tag;
  reg                 ways_0_metas_77_mru;
  reg                 ways_0_metas_78_vld;
  reg        [50:0]   ways_0_metas_78_tag;
  reg                 ways_0_metas_78_mru;
  reg                 ways_0_metas_79_vld;
  reg        [50:0]   ways_0_metas_79_tag;
  reg                 ways_0_metas_79_mru;
  reg                 ways_0_metas_80_vld;
  reg        [50:0]   ways_0_metas_80_tag;
  reg                 ways_0_metas_80_mru;
  reg                 ways_0_metas_81_vld;
  reg        [50:0]   ways_0_metas_81_tag;
  reg                 ways_0_metas_81_mru;
  reg                 ways_0_metas_82_vld;
  reg        [50:0]   ways_0_metas_82_tag;
  reg                 ways_0_metas_82_mru;
  reg                 ways_0_metas_83_vld;
  reg        [50:0]   ways_0_metas_83_tag;
  reg                 ways_0_metas_83_mru;
  reg                 ways_0_metas_84_vld;
  reg        [50:0]   ways_0_metas_84_tag;
  reg                 ways_0_metas_84_mru;
  reg                 ways_0_metas_85_vld;
  reg        [50:0]   ways_0_metas_85_tag;
  reg                 ways_0_metas_85_mru;
  reg                 ways_0_metas_86_vld;
  reg        [50:0]   ways_0_metas_86_tag;
  reg                 ways_0_metas_86_mru;
  reg                 ways_0_metas_87_vld;
  reg        [50:0]   ways_0_metas_87_tag;
  reg                 ways_0_metas_87_mru;
  reg                 ways_0_metas_88_vld;
  reg        [50:0]   ways_0_metas_88_tag;
  reg                 ways_0_metas_88_mru;
  reg                 ways_0_metas_89_vld;
  reg        [50:0]   ways_0_metas_89_tag;
  reg                 ways_0_metas_89_mru;
  reg                 ways_0_metas_90_vld;
  reg        [50:0]   ways_0_metas_90_tag;
  reg                 ways_0_metas_90_mru;
  reg                 ways_0_metas_91_vld;
  reg        [50:0]   ways_0_metas_91_tag;
  reg                 ways_0_metas_91_mru;
  reg                 ways_0_metas_92_vld;
  reg        [50:0]   ways_0_metas_92_tag;
  reg                 ways_0_metas_92_mru;
  reg                 ways_0_metas_93_vld;
  reg        [50:0]   ways_0_metas_93_tag;
  reg                 ways_0_metas_93_mru;
  reg                 ways_0_metas_94_vld;
  reg        [50:0]   ways_0_metas_94_tag;
  reg                 ways_0_metas_94_mru;
  reg                 ways_0_metas_95_vld;
  reg        [50:0]   ways_0_metas_95_tag;
  reg                 ways_0_metas_95_mru;
  reg                 ways_0_metas_96_vld;
  reg        [50:0]   ways_0_metas_96_tag;
  reg                 ways_0_metas_96_mru;
  reg                 ways_0_metas_97_vld;
  reg        [50:0]   ways_0_metas_97_tag;
  reg                 ways_0_metas_97_mru;
  reg                 ways_0_metas_98_vld;
  reg        [50:0]   ways_0_metas_98_tag;
  reg                 ways_0_metas_98_mru;
  reg                 ways_0_metas_99_vld;
  reg        [50:0]   ways_0_metas_99_tag;
  reg                 ways_0_metas_99_mru;
  reg                 ways_0_metas_100_vld;
  reg        [50:0]   ways_0_metas_100_tag;
  reg                 ways_0_metas_100_mru;
  reg                 ways_0_metas_101_vld;
  reg        [50:0]   ways_0_metas_101_tag;
  reg                 ways_0_metas_101_mru;
  reg                 ways_0_metas_102_vld;
  reg        [50:0]   ways_0_metas_102_tag;
  reg                 ways_0_metas_102_mru;
  reg                 ways_0_metas_103_vld;
  reg        [50:0]   ways_0_metas_103_tag;
  reg                 ways_0_metas_103_mru;
  reg                 ways_0_metas_104_vld;
  reg        [50:0]   ways_0_metas_104_tag;
  reg                 ways_0_metas_104_mru;
  reg                 ways_0_metas_105_vld;
  reg        [50:0]   ways_0_metas_105_tag;
  reg                 ways_0_metas_105_mru;
  reg                 ways_0_metas_106_vld;
  reg        [50:0]   ways_0_metas_106_tag;
  reg                 ways_0_metas_106_mru;
  reg                 ways_0_metas_107_vld;
  reg        [50:0]   ways_0_metas_107_tag;
  reg                 ways_0_metas_107_mru;
  reg                 ways_0_metas_108_vld;
  reg        [50:0]   ways_0_metas_108_tag;
  reg                 ways_0_metas_108_mru;
  reg                 ways_0_metas_109_vld;
  reg        [50:0]   ways_0_metas_109_tag;
  reg                 ways_0_metas_109_mru;
  reg                 ways_0_metas_110_vld;
  reg        [50:0]   ways_0_metas_110_tag;
  reg                 ways_0_metas_110_mru;
  reg                 ways_0_metas_111_vld;
  reg        [50:0]   ways_0_metas_111_tag;
  reg                 ways_0_metas_111_mru;
  reg                 ways_0_metas_112_vld;
  reg        [50:0]   ways_0_metas_112_tag;
  reg                 ways_0_metas_112_mru;
  reg                 ways_0_metas_113_vld;
  reg        [50:0]   ways_0_metas_113_tag;
  reg                 ways_0_metas_113_mru;
  reg                 ways_0_metas_114_vld;
  reg        [50:0]   ways_0_metas_114_tag;
  reg                 ways_0_metas_114_mru;
  reg                 ways_0_metas_115_vld;
  reg        [50:0]   ways_0_metas_115_tag;
  reg                 ways_0_metas_115_mru;
  reg                 ways_0_metas_116_vld;
  reg        [50:0]   ways_0_metas_116_tag;
  reg                 ways_0_metas_116_mru;
  reg                 ways_0_metas_117_vld;
  reg        [50:0]   ways_0_metas_117_tag;
  reg                 ways_0_metas_117_mru;
  reg                 ways_0_metas_118_vld;
  reg        [50:0]   ways_0_metas_118_tag;
  reg                 ways_0_metas_118_mru;
  reg                 ways_0_metas_119_vld;
  reg        [50:0]   ways_0_metas_119_tag;
  reg                 ways_0_metas_119_mru;
  reg                 ways_0_metas_120_vld;
  reg        [50:0]   ways_0_metas_120_tag;
  reg                 ways_0_metas_120_mru;
  reg                 ways_0_metas_121_vld;
  reg        [50:0]   ways_0_metas_121_tag;
  reg                 ways_0_metas_121_mru;
  reg                 ways_0_metas_122_vld;
  reg        [50:0]   ways_0_metas_122_tag;
  reg                 ways_0_metas_122_mru;
  reg                 ways_0_metas_123_vld;
  reg        [50:0]   ways_0_metas_123_tag;
  reg                 ways_0_metas_123_mru;
  reg                 ways_0_metas_124_vld;
  reg        [50:0]   ways_0_metas_124_tag;
  reg                 ways_0_metas_124_mru;
  reg                 ways_0_metas_125_vld;
  reg        [50:0]   ways_0_metas_125_tag;
  reg                 ways_0_metas_125_mru;
  reg                 ways_0_metas_126_vld;
  reg        [50:0]   ways_0_metas_126_tag;
  reg                 ways_0_metas_126_mru;
  reg                 ways_0_metas_127_vld;
  reg        [50:0]   ways_0_metas_127_tag;
  reg                 ways_0_metas_127_mru;
  reg                 ways_1_metas_0_vld;
  reg        [50:0]   ways_1_metas_0_tag;
  reg                 ways_1_metas_0_mru;
  reg                 ways_1_metas_1_vld;
  reg        [50:0]   ways_1_metas_1_tag;
  reg                 ways_1_metas_1_mru;
  reg                 ways_1_metas_2_vld;
  reg        [50:0]   ways_1_metas_2_tag;
  reg                 ways_1_metas_2_mru;
  reg                 ways_1_metas_3_vld;
  reg        [50:0]   ways_1_metas_3_tag;
  reg                 ways_1_metas_3_mru;
  reg                 ways_1_metas_4_vld;
  reg        [50:0]   ways_1_metas_4_tag;
  reg                 ways_1_metas_4_mru;
  reg                 ways_1_metas_5_vld;
  reg        [50:0]   ways_1_metas_5_tag;
  reg                 ways_1_metas_5_mru;
  reg                 ways_1_metas_6_vld;
  reg        [50:0]   ways_1_metas_6_tag;
  reg                 ways_1_metas_6_mru;
  reg                 ways_1_metas_7_vld;
  reg        [50:0]   ways_1_metas_7_tag;
  reg                 ways_1_metas_7_mru;
  reg                 ways_1_metas_8_vld;
  reg        [50:0]   ways_1_metas_8_tag;
  reg                 ways_1_metas_8_mru;
  reg                 ways_1_metas_9_vld;
  reg        [50:0]   ways_1_metas_9_tag;
  reg                 ways_1_metas_9_mru;
  reg                 ways_1_metas_10_vld;
  reg        [50:0]   ways_1_metas_10_tag;
  reg                 ways_1_metas_10_mru;
  reg                 ways_1_metas_11_vld;
  reg        [50:0]   ways_1_metas_11_tag;
  reg                 ways_1_metas_11_mru;
  reg                 ways_1_metas_12_vld;
  reg        [50:0]   ways_1_metas_12_tag;
  reg                 ways_1_metas_12_mru;
  reg                 ways_1_metas_13_vld;
  reg        [50:0]   ways_1_metas_13_tag;
  reg                 ways_1_metas_13_mru;
  reg                 ways_1_metas_14_vld;
  reg        [50:0]   ways_1_metas_14_tag;
  reg                 ways_1_metas_14_mru;
  reg                 ways_1_metas_15_vld;
  reg        [50:0]   ways_1_metas_15_tag;
  reg                 ways_1_metas_15_mru;
  reg                 ways_1_metas_16_vld;
  reg        [50:0]   ways_1_metas_16_tag;
  reg                 ways_1_metas_16_mru;
  reg                 ways_1_metas_17_vld;
  reg        [50:0]   ways_1_metas_17_tag;
  reg                 ways_1_metas_17_mru;
  reg                 ways_1_metas_18_vld;
  reg        [50:0]   ways_1_metas_18_tag;
  reg                 ways_1_metas_18_mru;
  reg                 ways_1_metas_19_vld;
  reg        [50:0]   ways_1_metas_19_tag;
  reg                 ways_1_metas_19_mru;
  reg                 ways_1_metas_20_vld;
  reg        [50:0]   ways_1_metas_20_tag;
  reg                 ways_1_metas_20_mru;
  reg                 ways_1_metas_21_vld;
  reg        [50:0]   ways_1_metas_21_tag;
  reg                 ways_1_metas_21_mru;
  reg                 ways_1_metas_22_vld;
  reg        [50:0]   ways_1_metas_22_tag;
  reg                 ways_1_metas_22_mru;
  reg                 ways_1_metas_23_vld;
  reg        [50:0]   ways_1_metas_23_tag;
  reg                 ways_1_metas_23_mru;
  reg                 ways_1_metas_24_vld;
  reg        [50:0]   ways_1_metas_24_tag;
  reg                 ways_1_metas_24_mru;
  reg                 ways_1_metas_25_vld;
  reg        [50:0]   ways_1_metas_25_tag;
  reg                 ways_1_metas_25_mru;
  reg                 ways_1_metas_26_vld;
  reg        [50:0]   ways_1_metas_26_tag;
  reg                 ways_1_metas_26_mru;
  reg                 ways_1_metas_27_vld;
  reg        [50:0]   ways_1_metas_27_tag;
  reg                 ways_1_metas_27_mru;
  reg                 ways_1_metas_28_vld;
  reg        [50:0]   ways_1_metas_28_tag;
  reg                 ways_1_metas_28_mru;
  reg                 ways_1_metas_29_vld;
  reg        [50:0]   ways_1_metas_29_tag;
  reg                 ways_1_metas_29_mru;
  reg                 ways_1_metas_30_vld;
  reg        [50:0]   ways_1_metas_30_tag;
  reg                 ways_1_metas_30_mru;
  reg                 ways_1_metas_31_vld;
  reg        [50:0]   ways_1_metas_31_tag;
  reg                 ways_1_metas_31_mru;
  reg                 ways_1_metas_32_vld;
  reg        [50:0]   ways_1_metas_32_tag;
  reg                 ways_1_metas_32_mru;
  reg                 ways_1_metas_33_vld;
  reg        [50:0]   ways_1_metas_33_tag;
  reg                 ways_1_metas_33_mru;
  reg                 ways_1_metas_34_vld;
  reg        [50:0]   ways_1_metas_34_tag;
  reg                 ways_1_metas_34_mru;
  reg                 ways_1_metas_35_vld;
  reg        [50:0]   ways_1_metas_35_tag;
  reg                 ways_1_metas_35_mru;
  reg                 ways_1_metas_36_vld;
  reg        [50:0]   ways_1_metas_36_tag;
  reg                 ways_1_metas_36_mru;
  reg                 ways_1_metas_37_vld;
  reg        [50:0]   ways_1_metas_37_tag;
  reg                 ways_1_metas_37_mru;
  reg                 ways_1_metas_38_vld;
  reg        [50:0]   ways_1_metas_38_tag;
  reg                 ways_1_metas_38_mru;
  reg                 ways_1_metas_39_vld;
  reg        [50:0]   ways_1_metas_39_tag;
  reg                 ways_1_metas_39_mru;
  reg                 ways_1_metas_40_vld;
  reg        [50:0]   ways_1_metas_40_tag;
  reg                 ways_1_metas_40_mru;
  reg                 ways_1_metas_41_vld;
  reg        [50:0]   ways_1_metas_41_tag;
  reg                 ways_1_metas_41_mru;
  reg                 ways_1_metas_42_vld;
  reg        [50:0]   ways_1_metas_42_tag;
  reg                 ways_1_metas_42_mru;
  reg                 ways_1_metas_43_vld;
  reg        [50:0]   ways_1_metas_43_tag;
  reg                 ways_1_metas_43_mru;
  reg                 ways_1_metas_44_vld;
  reg        [50:0]   ways_1_metas_44_tag;
  reg                 ways_1_metas_44_mru;
  reg                 ways_1_metas_45_vld;
  reg        [50:0]   ways_1_metas_45_tag;
  reg                 ways_1_metas_45_mru;
  reg                 ways_1_metas_46_vld;
  reg        [50:0]   ways_1_metas_46_tag;
  reg                 ways_1_metas_46_mru;
  reg                 ways_1_metas_47_vld;
  reg        [50:0]   ways_1_metas_47_tag;
  reg                 ways_1_metas_47_mru;
  reg                 ways_1_metas_48_vld;
  reg        [50:0]   ways_1_metas_48_tag;
  reg                 ways_1_metas_48_mru;
  reg                 ways_1_metas_49_vld;
  reg        [50:0]   ways_1_metas_49_tag;
  reg                 ways_1_metas_49_mru;
  reg                 ways_1_metas_50_vld;
  reg        [50:0]   ways_1_metas_50_tag;
  reg                 ways_1_metas_50_mru;
  reg                 ways_1_metas_51_vld;
  reg        [50:0]   ways_1_metas_51_tag;
  reg                 ways_1_metas_51_mru;
  reg                 ways_1_metas_52_vld;
  reg        [50:0]   ways_1_metas_52_tag;
  reg                 ways_1_metas_52_mru;
  reg                 ways_1_metas_53_vld;
  reg        [50:0]   ways_1_metas_53_tag;
  reg                 ways_1_metas_53_mru;
  reg                 ways_1_metas_54_vld;
  reg        [50:0]   ways_1_metas_54_tag;
  reg                 ways_1_metas_54_mru;
  reg                 ways_1_metas_55_vld;
  reg        [50:0]   ways_1_metas_55_tag;
  reg                 ways_1_metas_55_mru;
  reg                 ways_1_metas_56_vld;
  reg        [50:0]   ways_1_metas_56_tag;
  reg                 ways_1_metas_56_mru;
  reg                 ways_1_metas_57_vld;
  reg        [50:0]   ways_1_metas_57_tag;
  reg                 ways_1_metas_57_mru;
  reg                 ways_1_metas_58_vld;
  reg        [50:0]   ways_1_metas_58_tag;
  reg                 ways_1_metas_58_mru;
  reg                 ways_1_metas_59_vld;
  reg        [50:0]   ways_1_metas_59_tag;
  reg                 ways_1_metas_59_mru;
  reg                 ways_1_metas_60_vld;
  reg        [50:0]   ways_1_metas_60_tag;
  reg                 ways_1_metas_60_mru;
  reg                 ways_1_metas_61_vld;
  reg        [50:0]   ways_1_metas_61_tag;
  reg                 ways_1_metas_61_mru;
  reg                 ways_1_metas_62_vld;
  reg        [50:0]   ways_1_metas_62_tag;
  reg                 ways_1_metas_62_mru;
  reg                 ways_1_metas_63_vld;
  reg        [50:0]   ways_1_metas_63_tag;
  reg                 ways_1_metas_63_mru;
  reg                 ways_1_metas_64_vld;
  reg        [50:0]   ways_1_metas_64_tag;
  reg                 ways_1_metas_64_mru;
  reg                 ways_1_metas_65_vld;
  reg        [50:0]   ways_1_metas_65_tag;
  reg                 ways_1_metas_65_mru;
  reg                 ways_1_metas_66_vld;
  reg        [50:0]   ways_1_metas_66_tag;
  reg                 ways_1_metas_66_mru;
  reg                 ways_1_metas_67_vld;
  reg        [50:0]   ways_1_metas_67_tag;
  reg                 ways_1_metas_67_mru;
  reg                 ways_1_metas_68_vld;
  reg        [50:0]   ways_1_metas_68_tag;
  reg                 ways_1_metas_68_mru;
  reg                 ways_1_metas_69_vld;
  reg        [50:0]   ways_1_metas_69_tag;
  reg                 ways_1_metas_69_mru;
  reg                 ways_1_metas_70_vld;
  reg        [50:0]   ways_1_metas_70_tag;
  reg                 ways_1_metas_70_mru;
  reg                 ways_1_metas_71_vld;
  reg        [50:0]   ways_1_metas_71_tag;
  reg                 ways_1_metas_71_mru;
  reg                 ways_1_metas_72_vld;
  reg        [50:0]   ways_1_metas_72_tag;
  reg                 ways_1_metas_72_mru;
  reg                 ways_1_metas_73_vld;
  reg        [50:0]   ways_1_metas_73_tag;
  reg                 ways_1_metas_73_mru;
  reg                 ways_1_metas_74_vld;
  reg        [50:0]   ways_1_metas_74_tag;
  reg                 ways_1_metas_74_mru;
  reg                 ways_1_metas_75_vld;
  reg        [50:0]   ways_1_metas_75_tag;
  reg                 ways_1_metas_75_mru;
  reg                 ways_1_metas_76_vld;
  reg        [50:0]   ways_1_metas_76_tag;
  reg                 ways_1_metas_76_mru;
  reg                 ways_1_metas_77_vld;
  reg        [50:0]   ways_1_metas_77_tag;
  reg                 ways_1_metas_77_mru;
  reg                 ways_1_metas_78_vld;
  reg        [50:0]   ways_1_metas_78_tag;
  reg                 ways_1_metas_78_mru;
  reg                 ways_1_metas_79_vld;
  reg        [50:0]   ways_1_metas_79_tag;
  reg                 ways_1_metas_79_mru;
  reg                 ways_1_metas_80_vld;
  reg        [50:0]   ways_1_metas_80_tag;
  reg                 ways_1_metas_80_mru;
  reg                 ways_1_metas_81_vld;
  reg        [50:0]   ways_1_metas_81_tag;
  reg                 ways_1_metas_81_mru;
  reg                 ways_1_metas_82_vld;
  reg        [50:0]   ways_1_metas_82_tag;
  reg                 ways_1_metas_82_mru;
  reg                 ways_1_metas_83_vld;
  reg        [50:0]   ways_1_metas_83_tag;
  reg                 ways_1_metas_83_mru;
  reg                 ways_1_metas_84_vld;
  reg        [50:0]   ways_1_metas_84_tag;
  reg                 ways_1_metas_84_mru;
  reg                 ways_1_metas_85_vld;
  reg        [50:0]   ways_1_metas_85_tag;
  reg                 ways_1_metas_85_mru;
  reg                 ways_1_metas_86_vld;
  reg        [50:0]   ways_1_metas_86_tag;
  reg                 ways_1_metas_86_mru;
  reg                 ways_1_metas_87_vld;
  reg        [50:0]   ways_1_metas_87_tag;
  reg                 ways_1_metas_87_mru;
  reg                 ways_1_metas_88_vld;
  reg        [50:0]   ways_1_metas_88_tag;
  reg                 ways_1_metas_88_mru;
  reg                 ways_1_metas_89_vld;
  reg        [50:0]   ways_1_metas_89_tag;
  reg                 ways_1_metas_89_mru;
  reg                 ways_1_metas_90_vld;
  reg        [50:0]   ways_1_metas_90_tag;
  reg                 ways_1_metas_90_mru;
  reg                 ways_1_metas_91_vld;
  reg        [50:0]   ways_1_metas_91_tag;
  reg                 ways_1_metas_91_mru;
  reg                 ways_1_metas_92_vld;
  reg        [50:0]   ways_1_metas_92_tag;
  reg                 ways_1_metas_92_mru;
  reg                 ways_1_metas_93_vld;
  reg        [50:0]   ways_1_metas_93_tag;
  reg                 ways_1_metas_93_mru;
  reg                 ways_1_metas_94_vld;
  reg        [50:0]   ways_1_metas_94_tag;
  reg                 ways_1_metas_94_mru;
  reg                 ways_1_metas_95_vld;
  reg        [50:0]   ways_1_metas_95_tag;
  reg                 ways_1_metas_95_mru;
  reg                 ways_1_metas_96_vld;
  reg        [50:0]   ways_1_metas_96_tag;
  reg                 ways_1_metas_96_mru;
  reg                 ways_1_metas_97_vld;
  reg        [50:0]   ways_1_metas_97_tag;
  reg                 ways_1_metas_97_mru;
  reg                 ways_1_metas_98_vld;
  reg        [50:0]   ways_1_metas_98_tag;
  reg                 ways_1_metas_98_mru;
  reg                 ways_1_metas_99_vld;
  reg        [50:0]   ways_1_metas_99_tag;
  reg                 ways_1_metas_99_mru;
  reg                 ways_1_metas_100_vld;
  reg        [50:0]   ways_1_metas_100_tag;
  reg                 ways_1_metas_100_mru;
  reg                 ways_1_metas_101_vld;
  reg        [50:0]   ways_1_metas_101_tag;
  reg                 ways_1_metas_101_mru;
  reg                 ways_1_metas_102_vld;
  reg        [50:0]   ways_1_metas_102_tag;
  reg                 ways_1_metas_102_mru;
  reg                 ways_1_metas_103_vld;
  reg        [50:0]   ways_1_metas_103_tag;
  reg                 ways_1_metas_103_mru;
  reg                 ways_1_metas_104_vld;
  reg        [50:0]   ways_1_metas_104_tag;
  reg                 ways_1_metas_104_mru;
  reg                 ways_1_metas_105_vld;
  reg        [50:0]   ways_1_metas_105_tag;
  reg                 ways_1_metas_105_mru;
  reg                 ways_1_metas_106_vld;
  reg        [50:0]   ways_1_metas_106_tag;
  reg                 ways_1_metas_106_mru;
  reg                 ways_1_metas_107_vld;
  reg        [50:0]   ways_1_metas_107_tag;
  reg                 ways_1_metas_107_mru;
  reg                 ways_1_metas_108_vld;
  reg        [50:0]   ways_1_metas_108_tag;
  reg                 ways_1_metas_108_mru;
  reg                 ways_1_metas_109_vld;
  reg        [50:0]   ways_1_metas_109_tag;
  reg                 ways_1_metas_109_mru;
  reg                 ways_1_metas_110_vld;
  reg        [50:0]   ways_1_metas_110_tag;
  reg                 ways_1_metas_110_mru;
  reg                 ways_1_metas_111_vld;
  reg        [50:0]   ways_1_metas_111_tag;
  reg                 ways_1_metas_111_mru;
  reg                 ways_1_metas_112_vld;
  reg        [50:0]   ways_1_metas_112_tag;
  reg                 ways_1_metas_112_mru;
  reg                 ways_1_metas_113_vld;
  reg        [50:0]   ways_1_metas_113_tag;
  reg                 ways_1_metas_113_mru;
  reg                 ways_1_metas_114_vld;
  reg        [50:0]   ways_1_metas_114_tag;
  reg                 ways_1_metas_114_mru;
  reg                 ways_1_metas_115_vld;
  reg        [50:0]   ways_1_metas_115_tag;
  reg                 ways_1_metas_115_mru;
  reg                 ways_1_metas_116_vld;
  reg        [50:0]   ways_1_metas_116_tag;
  reg                 ways_1_metas_116_mru;
  reg                 ways_1_metas_117_vld;
  reg        [50:0]   ways_1_metas_117_tag;
  reg                 ways_1_metas_117_mru;
  reg                 ways_1_metas_118_vld;
  reg        [50:0]   ways_1_metas_118_tag;
  reg                 ways_1_metas_118_mru;
  reg                 ways_1_metas_119_vld;
  reg        [50:0]   ways_1_metas_119_tag;
  reg                 ways_1_metas_119_mru;
  reg                 ways_1_metas_120_vld;
  reg        [50:0]   ways_1_metas_120_tag;
  reg                 ways_1_metas_120_mru;
  reg                 ways_1_metas_121_vld;
  reg        [50:0]   ways_1_metas_121_tag;
  reg                 ways_1_metas_121_mru;
  reg                 ways_1_metas_122_vld;
  reg        [50:0]   ways_1_metas_122_tag;
  reg                 ways_1_metas_122_mru;
  reg                 ways_1_metas_123_vld;
  reg        [50:0]   ways_1_metas_123_tag;
  reg                 ways_1_metas_123_mru;
  reg                 ways_1_metas_124_vld;
  reg        [50:0]   ways_1_metas_124_tag;
  reg                 ways_1_metas_124_mru;
  reg                 ways_1_metas_125_vld;
  reg        [50:0]   ways_1_metas_125_tag;
  reg                 ways_1_metas_125_mru;
  reg                 ways_1_metas_126_vld;
  reg        [50:0]   ways_1_metas_126_tag;
  reg                 ways_1_metas_126_mru;
  reg                 ways_1_metas_127_vld;
  reg        [50:0]   ways_1_metas_127_tag;
  reg                 ways_1_metas_127_mru;
  reg                 ways_2_metas_0_vld;
  reg        [50:0]   ways_2_metas_0_tag;
  reg                 ways_2_metas_0_mru;
  reg                 ways_2_metas_1_vld;
  reg        [50:0]   ways_2_metas_1_tag;
  reg                 ways_2_metas_1_mru;
  reg                 ways_2_metas_2_vld;
  reg        [50:0]   ways_2_metas_2_tag;
  reg                 ways_2_metas_2_mru;
  reg                 ways_2_metas_3_vld;
  reg        [50:0]   ways_2_metas_3_tag;
  reg                 ways_2_metas_3_mru;
  reg                 ways_2_metas_4_vld;
  reg        [50:0]   ways_2_metas_4_tag;
  reg                 ways_2_metas_4_mru;
  reg                 ways_2_metas_5_vld;
  reg        [50:0]   ways_2_metas_5_tag;
  reg                 ways_2_metas_5_mru;
  reg                 ways_2_metas_6_vld;
  reg        [50:0]   ways_2_metas_6_tag;
  reg                 ways_2_metas_6_mru;
  reg                 ways_2_metas_7_vld;
  reg        [50:0]   ways_2_metas_7_tag;
  reg                 ways_2_metas_7_mru;
  reg                 ways_2_metas_8_vld;
  reg        [50:0]   ways_2_metas_8_tag;
  reg                 ways_2_metas_8_mru;
  reg                 ways_2_metas_9_vld;
  reg        [50:0]   ways_2_metas_9_tag;
  reg                 ways_2_metas_9_mru;
  reg                 ways_2_metas_10_vld;
  reg        [50:0]   ways_2_metas_10_tag;
  reg                 ways_2_metas_10_mru;
  reg                 ways_2_metas_11_vld;
  reg        [50:0]   ways_2_metas_11_tag;
  reg                 ways_2_metas_11_mru;
  reg                 ways_2_metas_12_vld;
  reg        [50:0]   ways_2_metas_12_tag;
  reg                 ways_2_metas_12_mru;
  reg                 ways_2_metas_13_vld;
  reg        [50:0]   ways_2_metas_13_tag;
  reg                 ways_2_metas_13_mru;
  reg                 ways_2_metas_14_vld;
  reg        [50:0]   ways_2_metas_14_tag;
  reg                 ways_2_metas_14_mru;
  reg                 ways_2_metas_15_vld;
  reg        [50:0]   ways_2_metas_15_tag;
  reg                 ways_2_metas_15_mru;
  reg                 ways_2_metas_16_vld;
  reg        [50:0]   ways_2_metas_16_tag;
  reg                 ways_2_metas_16_mru;
  reg                 ways_2_metas_17_vld;
  reg        [50:0]   ways_2_metas_17_tag;
  reg                 ways_2_metas_17_mru;
  reg                 ways_2_metas_18_vld;
  reg        [50:0]   ways_2_metas_18_tag;
  reg                 ways_2_metas_18_mru;
  reg                 ways_2_metas_19_vld;
  reg        [50:0]   ways_2_metas_19_tag;
  reg                 ways_2_metas_19_mru;
  reg                 ways_2_metas_20_vld;
  reg        [50:0]   ways_2_metas_20_tag;
  reg                 ways_2_metas_20_mru;
  reg                 ways_2_metas_21_vld;
  reg        [50:0]   ways_2_metas_21_tag;
  reg                 ways_2_metas_21_mru;
  reg                 ways_2_metas_22_vld;
  reg        [50:0]   ways_2_metas_22_tag;
  reg                 ways_2_metas_22_mru;
  reg                 ways_2_metas_23_vld;
  reg        [50:0]   ways_2_metas_23_tag;
  reg                 ways_2_metas_23_mru;
  reg                 ways_2_metas_24_vld;
  reg        [50:0]   ways_2_metas_24_tag;
  reg                 ways_2_metas_24_mru;
  reg                 ways_2_metas_25_vld;
  reg        [50:0]   ways_2_metas_25_tag;
  reg                 ways_2_metas_25_mru;
  reg                 ways_2_metas_26_vld;
  reg        [50:0]   ways_2_metas_26_tag;
  reg                 ways_2_metas_26_mru;
  reg                 ways_2_metas_27_vld;
  reg        [50:0]   ways_2_metas_27_tag;
  reg                 ways_2_metas_27_mru;
  reg                 ways_2_metas_28_vld;
  reg        [50:0]   ways_2_metas_28_tag;
  reg                 ways_2_metas_28_mru;
  reg                 ways_2_metas_29_vld;
  reg        [50:0]   ways_2_metas_29_tag;
  reg                 ways_2_metas_29_mru;
  reg                 ways_2_metas_30_vld;
  reg        [50:0]   ways_2_metas_30_tag;
  reg                 ways_2_metas_30_mru;
  reg                 ways_2_metas_31_vld;
  reg        [50:0]   ways_2_metas_31_tag;
  reg                 ways_2_metas_31_mru;
  reg                 ways_2_metas_32_vld;
  reg        [50:0]   ways_2_metas_32_tag;
  reg                 ways_2_metas_32_mru;
  reg                 ways_2_metas_33_vld;
  reg        [50:0]   ways_2_metas_33_tag;
  reg                 ways_2_metas_33_mru;
  reg                 ways_2_metas_34_vld;
  reg        [50:0]   ways_2_metas_34_tag;
  reg                 ways_2_metas_34_mru;
  reg                 ways_2_metas_35_vld;
  reg        [50:0]   ways_2_metas_35_tag;
  reg                 ways_2_metas_35_mru;
  reg                 ways_2_metas_36_vld;
  reg        [50:0]   ways_2_metas_36_tag;
  reg                 ways_2_metas_36_mru;
  reg                 ways_2_metas_37_vld;
  reg        [50:0]   ways_2_metas_37_tag;
  reg                 ways_2_metas_37_mru;
  reg                 ways_2_metas_38_vld;
  reg        [50:0]   ways_2_metas_38_tag;
  reg                 ways_2_metas_38_mru;
  reg                 ways_2_metas_39_vld;
  reg        [50:0]   ways_2_metas_39_tag;
  reg                 ways_2_metas_39_mru;
  reg                 ways_2_metas_40_vld;
  reg        [50:0]   ways_2_metas_40_tag;
  reg                 ways_2_metas_40_mru;
  reg                 ways_2_metas_41_vld;
  reg        [50:0]   ways_2_metas_41_tag;
  reg                 ways_2_metas_41_mru;
  reg                 ways_2_metas_42_vld;
  reg        [50:0]   ways_2_metas_42_tag;
  reg                 ways_2_metas_42_mru;
  reg                 ways_2_metas_43_vld;
  reg        [50:0]   ways_2_metas_43_tag;
  reg                 ways_2_metas_43_mru;
  reg                 ways_2_metas_44_vld;
  reg        [50:0]   ways_2_metas_44_tag;
  reg                 ways_2_metas_44_mru;
  reg                 ways_2_metas_45_vld;
  reg        [50:0]   ways_2_metas_45_tag;
  reg                 ways_2_metas_45_mru;
  reg                 ways_2_metas_46_vld;
  reg        [50:0]   ways_2_metas_46_tag;
  reg                 ways_2_metas_46_mru;
  reg                 ways_2_metas_47_vld;
  reg        [50:0]   ways_2_metas_47_tag;
  reg                 ways_2_metas_47_mru;
  reg                 ways_2_metas_48_vld;
  reg        [50:0]   ways_2_metas_48_tag;
  reg                 ways_2_metas_48_mru;
  reg                 ways_2_metas_49_vld;
  reg        [50:0]   ways_2_metas_49_tag;
  reg                 ways_2_metas_49_mru;
  reg                 ways_2_metas_50_vld;
  reg        [50:0]   ways_2_metas_50_tag;
  reg                 ways_2_metas_50_mru;
  reg                 ways_2_metas_51_vld;
  reg        [50:0]   ways_2_metas_51_tag;
  reg                 ways_2_metas_51_mru;
  reg                 ways_2_metas_52_vld;
  reg        [50:0]   ways_2_metas_52_tag;
  reg                 ways_2_metas_52_mru;
  reg                 ways_2_metas_53_vld;
  reg        [50:0]   ways_2_metas_53_tag;
  reg                 ways_2_metas_53_mru;
  reg                 ways_2_metas_54_vld;
  reg        [50:0]   ways_2_metas_54_tag;
  reg                 ways_2_metas_54_mru;
  reg                 ways_2_metas_55_vld;
  reg        [50:0]   ways_2_metas_55_tag;
  reg                 ways_2_metas_55_mru;
  reg                 ways_2_metas_56_vld;
  reg        [50:0]   ways_2_metas_56_tag;
  reg                 ways_2_metas_56_mru;
  reg                 ways_2_metas_57_vld;
  reg        [50:0]   ways_2_metas_57_tag;
  reg                 ways_2_metas_57_mru;
  reg                 ways_2_metas_58_vld;
  reg        [50:0]   ways_2_metas_58_tag;
  reg                 ways_2_metas_58_mru;
  reg                 ways_2_metas_59_vld;
  reg        [50:0]   ways_2_metas_59_tag;
  reg                 ways_2_metas_59_mru;
  reg                 ways_2_metas_60_vld;
  reg        [50:0]   ways_2_metas_60_tag;
  reg                 ways_2_metas_60_mru;
  reg                 ways_2_metas_61_vld;
  reg        [50:0]   ways_2_metas_61_tag;
  reg                 ways_2_metas_61_mru;
  reg                 ways_2_metas_62_vld;
  reg        [50:0]   ways_2_metas_62_tag;
  reg                 ways_2_metas_62_mru;
  reg                 ways_2_metas_63_vld;
  reg        [50:0]   ways_2_metas_63_tag;
  reg                 ways_2_metas_63_mru;
  reg                 ways_2_metas_64_vld;
  reg        [50:0]   ways_2_metas_64_tag;
  reg                 ways_2_metas_64_mru;
  reg                 ways_2_metas_65_vld;
  reg        [50:0]   ways_2_metas_65_tag;
  reg                 ways_2_metas_65_mru;
  reg                 ways_2_metas_66_vld;
  reg        [50:0]   ways_2_metas_66_tag;
  reg                 ways_2_metas_66_mru;
  reg                 ways_2_metas_67_vld;
  reg        [50:0]   ways_2_metas_67_tag;
  reg                 ways_2_metas_67_mru;
  reg                 ways_2_metas_68_vld;
  reg        [50:0]   ways_2_metas_68_tag;
  reg                 ways_2_metas_68_mru;
  reg                 ways_2_metas_69_vld;
  reg        [50:0]   ways_2_metas_69_tag;
  reg                 ways_2_metas_69_mru;
  reg                 ways_2_metas_70_vld;
  reg        [50:0]   ways_2_metas_70_tag;
  reg                 ways_2_metas_70_mru;
  reg                 ways_2_metas_71_vld;
  reg        [50:0]   ways_2_metas_71_tag;
  reg                 ways_2_metas_71_mru;
  reg                 ways_2_metas_72_vld;
  reg        [50:0]   ways_2_metas_72_tag;
  reg                 ways_2_metas_72_mru;
  reg                 ways_2_metas_73_vld;
  reg        [50:0]   ways_2_metas_73_tag;
  reg                 ways_2_metas_73_mru;
  reg                 ways_2_metas_74_vld;
  reg        [50:0]   ways_2_metas_74_tag;
  reg                 ways_2_metas_74_mru;
  reg                 ways_2_metas_75_vld;
  reg        [50:0]   ways_2_metas_75_tag;
  reg                 ways_2_metas_75_mru;
  reg                 ways_2_metas_76_vld;
  reg        [50:0]   ways_2_metas_76_tag;
  reg                 ways_2_metas_76_mru;
  reg                 ways_2_metas_77_vld;
  reg        [50:0]   ways_2_metas_77_tag;
  reg                 ways_2_metas_77_mru;
  reg                 ways_2_metas_78_vld;
  reg        [50:0]   ways_2_metas_78_tag;
  reg                 ways_2_metas_78_mru;
  reg                 ways_2_metas_79_vld;
  reg        [50:0]   ways_2_metas_79_tag;
  reg                 ways_2_metas_79_mru;
  reg                 ways_2_metas_80_vld;
  reg        [50:0]   ways_2_metas_80_tag;
  reg                 ways_2_metas_80_mru;
  reg                 ways_2_metas_81_vld;
  reg        [50:0]   ways_2_metas_81_tag;
  reg                 ways_2_metas_81_mru;
  reg                 ways_2_metas_82_vld;
  reg        [50:0]   ways_2_metas_82_tag;
  reg                 ways_2_metas_82_mru;
  reg                 ways_2_metas_83_vld;
  reg        [50:0]   ways_2_metas_83_tag;
  reg                 ways_2_metas_83_mru;
  reg                 ways_2_metas_84_vld;
  reg        [50:0]   ways_2_metas_84_tag;
  reg                 ways_2_metas_84_mru;
  reg                 ways_2_metas_85_vld;
  reg        [50:0]   ways_2_metas_85_tag;
  reg                 ways_2_metas_85_mru;
  reg                 ways_2_metas_86_vld;
  reg        [50:0]   ways_2_metas_86_tag;
  reg                 ways_2_metas_86_mru;
  reg                 ways_2_metas_87_vld;
  reg        [50:0]   ways_2_metas_87_tag;
  reg                 ways_2_metas_87_mru;
  reg                 ways_2_metas_88_vld;
  reg        [50:0]   ways_2_metas_88_tag;
  reg                 ways_2_metas_88_mru;
  reg                 ways_2_metas_89_vld;
  reg        [50:0]   ways_2_metas_89_tag;
  reg                 ways_2_metas_89_mru;
  reg                 ways_2_metas_90_vld;
  reg        [50:0]   ways_2_metas_90_tag;
  reg                 ways_2_metas_90_mru;
  reg                 ways_2_metas_91_vld;
  reg        [50:0]   ways_2_metas_91_tag;
  reg                 ways_2_metas_91_mru;
  reg                 ways_2_metas_92_vld;
  reg        [50:0]   ways_2_metas_92_tag;
  reg                 ways_2_metas_92_mru;
  reg                 ways_2_metas_93_vld;
  reg        [50:0]   ways_2_metas_93_tag;
  reg                 ways_2_metas_93_mru;
  reg                 ways_2_metas_94_vld;
  reg        [50:0]   ways_2_metas_94_tag;
  reg                 ways_2_metas_94_mru;
  reg                 ways_2_metas_95_vld;
  reg        [50:0]   ways_2_metas_95_tag;
  reg                 ways_2_metas_95_mru;
  reg                 ways_2_metas_96_vld;
  reg        [50:0]   ways_2_metas_96_tag;
  reg                 ways_2_metas_96_mru;
  reg                 ways_2_metas_97_vld;
  reg        [50:0]   ways_2_metas_97_tag;
  reg                 ways_2_metas_97_mru;
  reg                 ways_2_metas_98_vld;
  reg        [50:0]   ways_2_metas_98_tag;
  reg                 ways_2_metas_98_mru;
  reg                 ways_2_metas_99_vld;
  reg        [50:0]   ways_2_metas_99_tag;
  reg                 ways_2_metas_99_mru;
  reg                 ways_2_metas_100_vld;
  reg        [50:0]   ways_2_metas_100_tag;
  reg                 ways_2_metas_100_mru;
  reg                 ways_2_metas_101_vld;
  reg        [50:0]   ways_2_metas_101_tag;
  reg                 ways_2_metas_101_mru;
  reg                 ways_2_metas_102_vld;
  reg        [50:0]   ways_2_metas_102_tag;
  reg                 ways_2_metas_102_mru;
  reg                 ways_2_metas_103_vld;
  reg        [50:0]   ways_2_metas_103_tag;
  reg                 ways_2_metas_103_mru;
  reg                 ways_2_metas_104_vld;
  reg        [50:0]   ways_2_metas_104_tag;
  reg                 ways_2_metas_104_mru;
  reg                 ways_2_metas_105_vld;
  reg        [50:0]   ways_2_metas_105_tag;
  reg                 ways_2_metas_105_mru;
  reg                 ways_2_metas_106_vld;
  reg        [50:0]   ways_2_metas_106_tag;
  reg                 ways_2_metas_106_mru;
  reg                 ways_2_metas_107_vld;
  reg        [50:0]   ways_2_metas_107_tag;
  reg                 ways_2_metas_107_mru;
  reg                 ways_2_metas_108_vld;
  reg        [50:0]   ways_2_metas_108_tag;
  reg                 ways_2_metas_108_mru;
  reg                 ways_2_metas_109_vld;
  reg        [50:0]   ways_2_metas_109_tag;
  reg                 ways_2_metas_109_mru;
  reg                 ways_2_metas_110_vld;
  reg        [50:0]   ways_2_metas_110_tag;
  reg                 ways_2_metas_110_mru;
  reg                 ways_2_metas_111_vld;
  reg        [50:0]   ways_2_metas_111_tag;
  reg                 ways_2_metas_111_mru;
  reg                 ways_2_metas_112_vld;
  reg        [50:0]   ways_2_metas_112_tag;
  reg                 ways_2_metas_112_mru;
  reg                 ways_2_metas_113_vld;
  reg        [50:0]   ways_2_metas_113_tag;
  reg                 ways_2_metas_113_mru;
  reg                 ways_2_metas_114_vld;
  reg        [50:0]   ways_2_metas_114_tag;
  reg                 ways_2_metas_114_mru;
  reg                 ways_2_metas_115_vld;
  reg        [50:0]   ways_2_metas_115_tag;
  reg                 ways_2_metas_115_mru;
  reg                 ways_2_metas_116_vld;
  reg        [50:0]   ways_2_metas_116_tag;
  reg                 ways_2_metas_116_mru;
  reg                 ways_2_metas_117_vld;
  reg        [50:0]   ways_2_metas_117_tag;
  reg                 ways_2_metas_117_mru;
  reg                 ways_2_metas_118_vld;
  reg        [50:0]   ways_2_metas_118_tag;
  reg                 ways_2_metas_118_mru;
  reg                 ways_2_metas_119_vld;
  reg        [50:0]   ways_2_metas_119_tag;
  reg                 ways_2_metas_119_mru;
  reg                 ways_2_metas_120_vld;
  reg        [50:0]   ways_2_metas_120_tag;
  reg                 ways_2_metas_120_mru;
  reg                 ways_2_metas_121_vld;
  reg        [50:0]   ways_2_metas_121_tag;
  reg                 ways_2_metas_121_mru;
  reg                 ways_2_metas_122_vld;
  reg        [50:0]   ways_2_metas_122_tag;
  reg                 ways_2_metas_122_mru;
  reg                 ways_2_metas_123_vld;
  reg        [50:0]   ways_2_metas_123_tag;
  reg                 ways_2_metas_123_mru;
  reg                 ways_2_metas_124_vld;
  reg        [50:0]   ways_2_metas_124_tag;
  reg                 ways_2_metas_124_mru;
  reg                 ways_2_metas_125_vld;
  reg        [50:0]   ways_2_metas_125_tag;
  reg                 ways_2_metas_125_mru;
  reg                 ways_2_metas_126_vld;
  reg        [50:0]   ways_2_metas_126_tag;
  reg                 ways_2_metas_126_mru;
  reg                 ways_2_metas_127_vld;
  reg        [50:0]   ways_2_metas_127_tag;
  reg                 ways_2_metas_127_mru;
  reg                 ways_3_metas_0_vld;
  reg        [50:0]   ways_3_metas_0_tag;
  reg                 ways_3_metas_0_mru;
  reg                 ways_3_metas_1_vld;
  reg        [50:0]   ways_3_metas_1_tag;
  reg                 ways_3_metas_1_mru;
  reg                 ways_3_metas_2_vld;
  reg        [50:0]   ways_3_metas_2_tag;
  reg                 ways_3_metas_2_mru;
  reg                 ways_3_metas_3_vld;
  reg        [50:0]   ways_3_metas_3_tag;
  reg                 ways_3_metas_3_mru;
  reg                 ways_3_metas_4_vld;
  reg        [50:0]   ways_3_metas_4_tag;
  reg                 ways_3_metas_4_mru;
  reg                 ways_3_metas_5_vld;
  reg        [50:0]   ways_3_metas_5_tag;
  reg                 ways_3_metas_5_mru;
  reg                 ways_3_metas_6_vld;
  reg        [50:0]   ways_3_metas_6_tag;
  reg                 ways_3_metas_6_mru;
  reg                 ways_3_metas_7_vld;
  reg        [50:0]   ways_3_metas_7_tag;
  reg                 ways_3_metas_7_mru;
  reg                 ways_3_metas_8_vld;
  reg        [50:0]   ways_3_metas_8_tag;
  reg                 ways_3_metas_8_mru;
  reg                 ways_3_metas_9_vld;
  reg        [50:0]   ways_3_metas_9_tag;
  reg                 ways_3_metas_9_mru;
  reg                 ways_3_metas_10_vld;
  reg        [50:0]   ways_3_metas_10_tag;
  reg                 ways_3_metas_10_mru;
  reg                 ways_3_metas_11_vld;
  reg        [50:0]   ways_3_metas_11_tag;
  reg                 ways_3_metas_11_mru;
  reg                 ways_3_metas_12_vld;
  reg        [50:0]   ways_3_metas_12_tag;
  reg                 ways_3_metas_12_mru;
  reg                 ways_3_metas_13_vld;
  reg        [50:0]   ways_3_metas_13_tag;
  reg                 ways_3_metas_13_mru;
  reg                 ways_3_metas_14_vld;
  reg        [50:0]   ways_3_metas_14_tag;
  reg                 ways_3_metas_14_mru;
  reg                 ways_3_metas_15_vld;
  reg        [50:0]   ways_3_metas_15_tag;
  reg                 ways_3_metas_15_mru;
  reg                 ways_3_metas_16_vld;
  reg        [50:0]   ways_3_metas_16_tag;
  reg                 ways_3_metas_16_mru;
  reg                 ways_3_metas_17_vld;
  reg        [50:0]   ways_3_metas_17_tag;
  reg                 ways_3_metas_17_mru;
  reg                 ways_3_metas_18_vld;
  reg        [50:0]   ways_3_metas_18_tag;
  reg                 ways_3_metas_18_mru;
  reg                 ways_3_metas_19_vld;
  reg        [50:0]   ways_3_metas_19_tag;
  reg                 ways_3_metas_19_mru;
  reg                 ways_3_metas_20_vld;
  reg        [50:0]   ways_3_metas_20_tag;
  reg                 ways_3_metas_20_mru;
  reg                 ways_3_metas_21_vld;
  reg        [50:0]   ways_3_metas_21_tag;
  reg                 ways_3_metas_21_mru;
  reg                 ways_3_metas_22_vld;
  reg        [50:0]   ways_3_metas_22_tag;
  reg                 ways_3_metas_22_mru;
  reg                 ways_3_metas_23_vld;
  reg        [50:0]   ways_3_metas_23_tag;
  reg                 ways_3_metas_23_mru;
  reg                 ways_3_metas_24_vld;
  reg        [50:0]   ways_3_metas_24_tag;
  reg                 ways_3_metas_24_mru;
  reg                 ways_3_metas_25_vld;
  reg        [50:0]   ways_3_metas_25_tag;
  reg                 ways_3_metas_25_mru;
  reg                 ways_3_metas_26_vld;
  reg        [50:0]   ways_3_metas_26_tag;
  reg                 ways_3_metas_26_mru;
  reg                 ways_3_metas_27_vld;
  reg        [50:0]   ways_3_metas_27_tag;
  reg                 ways_3_metas_27_mru;
  reg                 ways_3_metas_28_vld;
  reg        [50:0]   ways_3_metas_28_tag;
  reg                 ways_3_metas_28_mru;
  reg                 ways_3_metas_29_vld;
  reg        [50:0]   ways_3_metas_29_tag;
  reg                 ways_3_metas_29_mru;
  reg                 ways_3_metas_30_vld;
  reg        [50:0]   ways_3_metas_30_tag;
  reg                 ways_3_metas_30_mru;
  reg                 ways_3_metas_31_vld;
  reg        [50:0]   ways_3_metas_31_tag;
  reg                 ways_3_metas_31_mru;
  reg                 ways_3_metas_32_vld;
  reg        [50:0]   ways_3_metas_32_tag;
  reg                 ways_3_metas_32_mru;
  reg                 ways_3_metas_33_vld;
  reg        [50:0]   ways_3_metas_33_tag;
  reg                 ways_3_metas_33_mru;
  reg                 ways_3_metas_34_vld;
  reg        [50:0]   ways_3_metas_34_tag;
  reg                 ways_3_metas_34_mru;
  reg                 ways_3_metas_35_vld;
  reg        [50:0]   ways_3_metas_35_tag;
  reg                 ways_3_metas_35_mru;
  reg                 ways_3_metas_36_vld;
  reg        [50:0]   ways_3_metas_36_tag;
  reg                 ways_3_metas_36_mru;
  reg                 ways_3_metas_37_vld;
  reg        [50:0]   ways_3_metas_37_tag;
  reg                 ways_3_metas_37_mru;
  reg                 ways_3_metas_38_vld;
  reg        [50:0]   ways_3_metas_38_tag;
  reg                 ways_3_metas_38_mru;
  reg                 ways_3_metas_39_vld;
  reg        [50:0]   ways_3_metas_39_tag;
  reg                 ways_3_metas_39_mru;
  reg                 ways_3_metas_40_vld;
  reg        [50:0]   ways_3_metas_40_tag;
  reg                 ways_3_metas_40_mru;
  reg                 ways_3_metas_41_vld;
  reg        [50:0]   ways_3_metas_41_tag;
  reg                 ways_3_metas_41_mru;
  reg                 ways_3_metas_42_vld;
  reg        [50:0]   ways_3_metas_42_tag;
  reg                 ways_3_metas_42_mru;
  reg                 ways_3_metas_43_vld;
  reg        [50:0]   ways_3_metas_43_tag;
  reg                 ways_3_metas_43_mru;
  reg                 ways_3_metas_44_vld;
  reg        [50:0]   ways_3_metas_44_tag;
  reg                 ways_3_metas_44_mru;
  reg                 ways_3_metas_45_vld;
  reg        [50:0]   ways_3_metas_45_tag;
  reg                 ways_3_metas_45_mru;
  reg                 ways_3_metas_46_vld;
  reg        [50:0]   ways_3_metas_46_tag;
  reg                 ways_3_metas_46_mru;
  reg                 ways_3_metas_47_vld;
  reg        [50:0]   ways_3_metas_47_tag;
  reg                 ways_3_metas_47_mru;
  reg                 ways_3_metas_48_vld;
  reg        [50:0]   ways_3_metas_48_tag;
  reg                 ways_3_metas_48_mru;
  reg                 ways_3_metas_49_vld;
  reg        [50:0]   ways_3_metas_49_tag;
  reg                 ways_3_metas_49_mru;
  reg                 ways_3_metas_50_vld;
  reg        [50:0]   ways_3_metas_50_tag;
  reg                 ways_3_metas_50_mru;
  reg                 ways_3_metas_51_vld;
  reg        [50:0]   ways_3_metas_51_tag;
  reg                 ways_3_metas_51_mru;
  reg                 ways_3_metas_52_vld;
  reg        [50:0]   ways_3_metas_52_tag;
  reg                 ways_3_metas_52_mru;
  reg                 ways_3_metas_53_vld;
  reg        [50:0]   ways_3_metas_53_tag;
  reg                 ways_3_metas_53_mru;
  reg                 ways_3_metas_54_vld;
  reg        [50:0]   ways_3_metas_54_tag;
  reg                 ways_3_metas_54_mru;
  reg                 ways_3_metas_55_vld;
  reg        [50:0]   ways_3_metas_55_tag;
  reg                 ways_3_metas_55_mru;
  reg                 ways_3_metas_56_vld;
  reg        [50:0]   ways_3_metas_56_tag;
  reg                 ways_3_metas_56_mru;
  reg                 ways_3_metas_57_vld;
  reg        [50:0]   ways_3_metas_57_tag;
  reg                 ways_3_metas_57_mru;
  reg                 ways_3_metas_58_vld;
  reg        [50:0]   ways_3_metas_58_tag;
  reg                 ways_3_metas_58_mru;
  reg                 ways_3_metas_59_vld;
  reg        [50:0]   ways_3_metas_59_tag;
  reg                 ways_3_metas_59_mru;
  reg                 ways_3_metas_60_vld;
  reg        [50:0]   ways_3_metas_60_tag;
  reg                 ways_3_metas_60_mru;
  reg                 ways_3_metas_61_vld;
  reg        [50:0]   ways_3_metas_61_tag;
  reg                 ways_3_metas_61_mru;
  reg                 ways_3_metas_62_vld;
  reg        [50:0]   ways_3_metas_62_tag;
  reg                 ways_3_metas_62_mru;
  reg                 ways_3_metas_63_vld;
  reg        [50:0]   ways_3_metas_63_tag;
  reg                 ways_3_metas_63_mru;
  reg                 ways_3_metas_64_vld;
  reg        [50:0]   ways_3_metas_64_tag;
  reg                 ways_3_metas_64_mru;
  reg                 ways_3_metas_65_vld;
  reg        [50:0]   ways_3_metas_65_tag;
  reg                 ways_3_metas_65_mru;
  reg                 ways_3_metas_66_vld;
  reg        [50:0]   ways_3_metas_66_tag;
  reg                 ways_3_metas_66_mru;
  reg                 ways_3_metas_67_vld;
  reg        [50:0]   ways_3_metas_67_tag;
  reg                 ways_3_metas_67_mru;
  reg                 ways_3_metas_68_vld;
  reg        [50:0]   ways_3_metas_68_tag;
  reg                 ways_3_metas_68_mru;
  reg                 ways_3_metas_69_vld;
  reg        [50:0]   ways_3_metas_69_tag;
  reg                 ways_3_metas_69_mru;
  reg                 ways_3_metas_70_vld;
  reg        [50:0]   ways_3_metas_70_tag;
  reg                 ways_3_metas_70_mru;
  reg                 ways_3_metas_71_vld;
  reg        [50:0]   ways_3_metas_71_tag;
  reg                 ways_3_metas_71_mru;
  reg                 ways_3_metas_72_vld;
  reg        [50:0]   ways_3_metas_72_tag;
  reg                 ways_3_metas_72_mru;
  reg                 ways_3_metas_73_vld;
  reg        [50:0]   ways_3_metas_73_tag;
  reg                 ways_3_metas_73_mru;
  reg                 ways_3_metas_74_vld;
  reg        [50:0]   ways_3_metas_74_tag;
  reg                 ways_3_metas_74_mru;
  reg                 ways_3_metas_75_vld;
  reg        [50:0]   ways_3_metas_75_tag;
  reg                 ways_3_metas_75_mru;
  reg                 ways_3_metas_76_vld;
  reg        [50:0]   ways_3_metas_76_tag;
  reg                 ways_3_metas_76_mru;
  reg                 ways_3_metas_77_vld;
  reg        [50:0]   ways_3_metas_77_tag;
  reg                 ways_3_metas_77_mru;
  reg                 ways_3_metas_78_vld;
  reg        [50:0]   ways_3_metas_78_tag;
  reg                 ways_3_metas_78_mru;
  reg                 ways_3_metas_79_vld;
  reg        [50:0]   ways_3_metas_79_tag;
  reg                 ways_3_metas_79_mru;
  reg                 ways_3_metas_80_vld;
  reg        [50:0]   ways_3_metas_80_tag;
  reg                 ways_3_metas_80_mru;
  reg                 ways_3_metas_81_vld;
  reg        [50:0]   ways_3_metas_81_tag;
  reg                 ways_3_metas_81_mru;
  reg                 ways_3_metas_82_vld;
  reg        [50:0]   ways_3_metas_82_tag;
  reg                 ways_3_metas_82_mru;
  reg                 ways_3_metas_83_vld;
  reg        [50:0]   ways_3_metas_83_tag;
  reg                 ways_3_metas_83_mru;
  reg                 ways_3_metas_84_vld;
  reg        [50:0]   ways_3_metas_84_tag;
  reg                 ways_3_metas_84_mru;
  reg                 ways_3_metas_85_vld;
  reg        [50:0]   ways_3_metas_85_tag;
  reg                 ways_3_metas_85_mru;
  reg                 ways_3_metas_86_vld;
  reg        [50:0]   ways_3_metas_86_tag;
  reg                 ways_3_metas_86_mru;
  reg                 ways_3_metas_87_vld;
  reg        [50:0]   ways_3_metas_87_tag;
  reg                 ways_3_metas_87_mru;
  reg                 ways_3_metas_88_vld;
  reg        [50:0]   ways_3_metas_88_tag;
  reg                 ways_3_metas_88_mru;
  reg                 ways_3_metas_89_vld;
  reg        [50:0]   ways_3_metas_89_tag;
  reg                 ways_3_metas_89_mru;
  reg                 ways_3_metas_90_vld;
  reg        [50:0]   ways_3_metas_90_tag;
  reg                 ways_3_metas_90_mru;
  reg                 ways_3_metas_91_vld;
  reg        [50:0]   ways_3_metas_91_tag;
  reg                 ways_3_metas_91_mru;
  reg                 ways_3_metas_92_vld;
  reg        [50:0]   ways_3_metas_92_tag;
  reg                 ways_3_metas_92_mru;
  reg                 ways_3_metas_93_vld;
  reg        [50:0]   ways_3_metas_93_tag;
  reg                 ways_3_metas_93_mru;
  reg                 ways_3_metas_94_vld;
  reg        [50:0]   ways_3_metas_94_tag;
  reg                 ways_3_metas_94_mru;
  reg                 ways_3_metas_95_vld;
  reg        [50:0]   ways_3_metas_95_tag;
  reg                 ways_3_metas_95_mru;
  reg                 ways_3_metas_96_vld;
  reg        [50:0]   ways_3_metas_96_tag;
  reg                 ways_3_metas_96_mru;
  reg                 ways_3_metas_97_vld;
  reg        [50:0]   ways_3_metas_97_tag;
  reg                 ways_3_metas_97_mru;
  reg                 ways_3_metas_98_vld;
  reg        [50:0]   ways_3_metas_98_tag;
  reg                 ways_3_metas_98_mru;
  reg                 ways_3_metas_99_vld;
  reg        [50:0]   ways_3_metas_99_tag;
  reg                 ways_3_metas_99_mru;
  reg                 ways_3_metas_100_vld;
  reg        [50:0]   ways_3_metas_100_tag;
  reg                 ways_3_metas_100_mru;
  reg                 ways_3_metas_101_vld;
  reg        [50:0]   ways_3_metas_101_tag;
  reg                 ways_3_metas_101_mru;
  reg                 ways_3_metas_102_vld;
  reg        [50:0]   ways_3_metas_102_tag;
  reg                 ways_3_metas_102_mru;
  reg                 ways_3_metas_103_vld;
  reg        [50:0]   ways_3_metas_103_tag;
  reg                 ways_3_metas_103_mru;
  reg                 ways_3_metas_104_vld;
  reg        [50:0]   ways_3_metas_104_tag;
  reg                 ways_3_metas_104_mru;
  reg                 ways_3_metas_105_vld;
  reg        [50:0]   ways_3_metas_105_tag;
  reg                 ways_3_metas_105_mru;
  reg                 ways_3_metas_106_vld;
  reg        [50:0]   ways_3_metas_106_tag;
  reg                 ways_3_metas_106_mru;
  reg                 ways_3_metas_107_vld;
  reg        [50:0]   ways_3_metas_107_tag;
  reg                 ways_3_metas_107_mru;
  reg                 ways_3_metas_108_vld;
  reg        [50:0]   ways_3_metas_108_tag;
  reg                 ways_3_metas_108_mru;
  reg                 ways_3_metas_109_vld;
  reg        [50:0]   ways_3_metas_109_tag;
  reg                 ways_3_metas_109_mru;
  reg                 ways_3_metas_110_vld;
  reg        [50:0]   ways_3_metas_110_tag;
  reg                 ways_3_metas_110_mru;
  reg                 ways_3_metas_111_vld;
  reg        [50:0]   ways_3_metas_111_tag;
  reg                 ways_3_metas_111_mru;
  reg                 ways_3_metas_112_vld;
  reg        [50:0]   ways_3_metas_112_tag;
  reg                 ways_3_metas_112_mru;
  reg                 ways_3_metas_113_vld;
  reg        [50:0]   ways_3_metas_113_tag;
  reg                 ways_3_metas_113_mru;
  reg                 ways_3_metas_114_vld;
  reg        [50:0]   ways_3_metas_114_tag;
  reg                 ways_3_metas_114_mru;
  reg                 ways_3_metas_115_vld;
  reg        [50:0]   ways_3_metas_115_tag;
  reg                 ways_3_metas_115_mru;
  reg                 ways_3_metas_116_vld;
  reg        [50:0]   ways_3_metas_116_tag;
  reg                 ways_3_metas_116_mru;
  reg                 ways_3_metas_117_vld;
  reg        [50:0]   ways_3_metas_117_tag;
  reg                 ways_3_metas_117_mru;
  reg                 ways_3_metas_118_vld;
  reg        [50:0]   ways_3_metas_118_tag;
  reg                 ways_3_metas_118_mru;
  reg                 ways_3_metas_119_vld;
  reg        [50:0]   ways_3_metas_119_tag;
  reg                 ways_3_metas_119_mru;
  reg                 ways_3_metas_120_vld;
  reg        [50:0]   ways_3_metas_120_tag;
  reg                 ways_3_metas_120_mru;
  reg                 ways_3_metas_121_vld;
  reg        [50:0]   ways_3_metas_121_tag;
  reg                 ways_3_metas_121_mru;
  reg                 ways_3_metas_122_vld;
  reg        [50:0]   ways_3_metas_122_tag;
  reg                 ways_3_metas_122_mru;
  reg                 ways_3_metas_123_vld;
  reg        [50:0]   ways_3_metas_123_tag;
  reg                 ways_3_metas_123_mru;
  reg                 ways_3_metas_124_vld;
  reg        [50:0]   ways_3_metas_124_tag;
  reg                 ways_3_metas_124_mru;
  reg                 ways_3_metas_125_vld;
  reg        [50:0]   ways_3_metas_125_tag;
  reg                 ways_3_metas_125_mru;
  reg                 ways_3_metas_126_vld;
  reg        [50:0]   ways_3_metas_126_tag;
  reg                 ways_3_metas_126_mru;
  reg                 ways_3_metas_127_vld;
  reg        [50:0]   ways_3_metas_127_tag;
  reg                 ways_3_metas_127_mru;
  wire       [50:0]   cache_tag_0;
  wire       [50:0]   cache_tag_1;
  wire       [50:0]   cache_tag_2;
  wire       [50:0]   cache_tag_3;
  wire                cache_hit_0;
  wire                cache_hit_1;
  wire                cache_hit_2;
  wire                cache_hit_3;
  wire                cache_invld_0;
  wire                cache_invld_1;
  wire                cache_invld_2;
  wire                cache_invld_3;
  wire                cache_victim_0;
  wire                cache_victim_1;
  wire                cache_victim_2;
  wire                cache_victim_3;
  wire                cache_mru_0;
  wire                cache_mru_1;
  wire                cache_mru_2;
  wire                cache_mru_3;
  wire                cache_lru_0;
  wire                cache_lru_1;
  wire                cache_lru_2;
  wire                cache_lru_3;
  wire       [1:0]    hit_id;
  wire       [1:0]    evict_id;
  wire       [1:0]    invld_id;
  wire       [1:0]    victim_id;
  wire                mru_full;
  wire                cpu_cmd_fire;
  wire                is_hit;
  wire                cpu_cmd_fire_1;
  wire                is_miss;
  wire                is_diff;
  wire                cpu_cmd_fire_2;
  wire                is_write;
  reg                 flush_busy;
  reg                 flush_cnt_willIncrement;
  reg                 flush_cnt_willClear;
  reg        [6:0]    flush_cnt_valueNext;
  reg        [6:0]    flush_cnt_value;
  wire                flush_cnt_willOverflowIfInc;
  wire                flush_cnt_willOverflow;
  wire                flush_done;
  wire                cache_hit_gnt_0;
  wire                cache_hit_gnt_1;
  wire                cache_hit_gnt_2;
  wire                cache_hit_gnt_3;
  wire                cache_victim_gnt_0;
  wire                cache_victim_gnt_1;
  wire                cache_victim_gnt_2;
  wire                cache_victim_gnt_3;
  wire                cache_invld_gnt_0;
  wire                cache_invld_gnt_1;
  wire                cache_invld_gnt_2;
  wire                cache_invld_gnt_3;
  reg        [1:0]    evict_id_miss;
  reg                 cpu_cmd_ready_1;
  wire       [50:0]   cpu_tag;
  wire       [6:0]    cpu_set;
  wire       [6:0]    cpu_bank_addr;
  wire       [2:0]    cpu_bank_index;
  wire       [511:0]  sram_banks_data_0;
  wire       [511:0]  sram_banks_data_1;
  wire       [511:0]  sram_banks_data_2;
  wire       [511:0]  sram_banks_data_3;
  wire                sram_banks_valid_0;
  wire                sram_banks_valid_1;
  wire                sram_banks_valid_2;
  wire                sram_banks_valid_3;
  reg                 next_level_cmd_valid_1;
  reg                 next_level_data_cnt_willIncrement;
  reg                 next_level_data_cnt_willClear;
  reg        [2:0]    next_level_data_cnt_valueNext;
  reg        [2:0]    next_level_data_cnt_value;
  wire                next_level_data_cnt_willOverflowIfInc;
  wire                next_level_data_cnt_willOverflow;
  wire       [6:0]    next_level_bank_addr;
  wire                next_level_rvalid;
  reg                 next_level_rdone;
  reg                 next_level_wdone;
  wire       [7:0]    next_level_wstrb_tmp;
  wire       [63:0]   next_level_wdata_tmp;
  wire       [7:0]    next_level_wstrb;
  wire       [63:0]   next_level_wdata;
  wire                when_DCache_l123;
  wire                when_DCache_l131;
  wire                when_DCache_l149;
  wire       [3:0]    _zz_cache_hit_gnt_0;
  wire       [3:0]    _zz_cache_hit_gnt_0_1;
  wire       [7:0]    _zz_cache_hit_gnt_0_2;
  wire       [7:0]    _zz_cache_hit_gnt_0_3;
  wire       [3:0]    _zz_cache_hit_gnt_0_4;
  wire       [3:0]    _zz_cache_invld_gnt_0;
  wire       [3:0]    _zz_cache_invld_gnt_0_1;
  wire       [7:0]    _zz_cache_invld_gnt_0_2;
  wire       [7:0]    _zz_cache_invld_gnt_0_3;
  wire       [3:0]    _zz_cache_invld_gnt_0_4;
  wire       [3:0]    _zz_cache_victim_gnt_0;
  wire       [3:0]    _zz_cache_victim_gnt_0_1;
  wire       [7:0]    _zz_cache_victim_gnt_0_2;
  wire       [7:0]    _zz_cache_victim_gnt_0_3;
  wire       [3:0]    _zz_cache_victim_gnt_0_4;
  wire                _zz_hit_id;
  wire                _zz_hit_id_1;
  wire                _zz_invld_id;
  wire                _zz_invld_id_1;
  wire                _zz_victim_id;
  wire                _zz_victim_id_1;
  wire                _zz_cache_hit_0;
  wire                _zz_cache_mru_0;
  wire       [127:0]  _zz_1;
  wire                _zz_2;
  wire                _zz_3;
  wire                _zz_4;
  wire                _zz_5;
  wire                _zz_6;
  wire                _zz_7;
  wire                _zz_8;
  wire                _zz_9;
  wire                _zz_10;
  wire                _zz_11;
  wire                _zz_12;
  wire                _zz_13;
  wire                _zz_14;
  wire                _zz_15;
  wire                _zz_16;
  wire                _zz_17;
  wire                _zz_18;
  wire                _zz_19;
  wire                _zz_20;
  wire                _zz_21;
  wire                _zz_22;
  wire                _zz_23;
  wire                _zz_24;
  wire                _zz_25;
  wire                _zz_26;
  wire                _zz_27;
  wire                _zz_28;
  wire                _zz_29;
  wire                _zz_30;
  wire                _zz_31;
  wire                _zz_32;
  wire                _zz_33;
  wire                _zz_34;
  wire                _zz_35;
  wire                _zz_36;
  wire                _zz_37;
  wire                _zz_38;
  wire                _zz_39;
  wire                _zz_40;
  wire                _zz_41;
  wire                _zz_42;
  wire                _zz_43;
  wire                _zz_44;
  wire                _zz_45;
  wire                _zz_46;
  wire                _zz_47;
  wire                _zz_48;
  wire                _zz_49;
  wire                _zz_50;
  wire                _zz_51;
  wire                _zz_52;
  wire                _zz_53;
  wire                _zz_54;
  wire                _zz_55;
  wire                _zz_56;
  wire                _zz_57;
  wire                _zz_58;
  wire                _zz_59;
  wire                _zz_60;
  wire                _zz_61;
  wire                _zz_62;
  wire                _zz_63;
  wire                _zz_64;
  wire                _zz_65;
  wire                _zz_66;
  wire                _zz_67;
  wire                _zz_68;
  wire                _zz_69;
  wire                _zz_70;
  wire                _zz_71;
  wire                _zz_72;
  wire                _zz_73;
  wire                _zz_74;
  wire                _zz_75;
  wire                _zz_76;
  wire                _zz_77;
  wire                _zz_78;
  wire                _zz_79;
  wire                _zz_80;
  wire                _zz_81;
  wire                _zz_82;
  wire                _zz_83;
  wire                _zz_84;
  wire                _zz_85;
  wire                _zz_86;
  wire                _zz_87;
  wire                _zz_88;
  wire                _zz_89;
  wire                _zz_90;
  wire                _zz_91;
  wire                _zz_92;
  wire                _zz_93;
  wire                _zz_94;
  wire                _zz_95;
  wire                _zz_96;
  wire                _zz_97;
  wire                _zz_98;
  wire                _zz_99;
  wire                _zz_100;
  wire                _zz_101;
  wire                _zz_102;
  wire                _zz_103;
  wire                _zz_104;
  wire                _zz_105;
  wire                _zz_106;
  wire                _zz_107;
  wire                _zz_108;
  wire                _zz_109;
  wire                _zz_110;
  wire                _zz_111;
  wire                _zz_112;
  wire                _zz_113;
  wire                _zz_114;
  wire                _zz_115;
  wire                _zz_116;
  wire                _zz_117;
  wire                _zz_118;
  wire                _zz_119;
  wire                _zz_120;
  wire                _zz_121;
  wire                _zz_122;
  wire                _zz_123;
  wire                _zz_124;
  wire                _zz_125;
  wire                _zz_126;
  wire                _zz_127;
  wire                _zz_128;
  wire                _zz_129;
  wire                when_DCache_l181;
  reg        [7:0]    _zz_sram_0_ports_cmd_payload_wen;
  wire                when_DCache_l188;
  wire                when_DCache_l195;
  wire       [127:0]  _zz_130;
  wire                _zz_131;
  wire                _zz_132;
  wire                _zz_133;
  wire                _zz_134;
  wire                _zz_135;
  wire                _zz_136;
  wire                _zz_137;
  wire                _zz_138;
  wire                _zz_139;
  wire                _zz_140;
  wire                _zz_141;
  wire                _zz_142;
  wire                _zz_143;
  wire                _zz_144;
  wire                _zz_145;
  wire                _zz_146;
  wire                _zz_147;
  wire                _zz_148;
  wire                _zz_149;
  wire                _zz_150;
  wire                _zz_151;
  wire                _zz_152;
  wire                _zz_153;
  wire                _zz_154;
  wire                _zz_155;
  wire                _zz_156;
  wire                _zz_157;
  wire                _zz_158;
  wire                _zz_159;
  wire                _zz_160;
  wire                _zz_161;
  wire                _zz_162;
  wire                _zz_163;
  wire                _zz_164;
  wire                _zz_165;
  wire                _zz_166;
  wire                _zz_167;
  wire                _zz_168;
  wire                _zz_169;
  wire                _zz_170;
  wire                _zz_171;
  wire                _zz_172;
  wire                _zz_173;
  wire                _zz_174;
  wire                _zz_175;
  wire                _zz_176;
  wire                _zz_177;
  wire                _zz_178;
  wire                _zz_179;
  wire                _zz_180;
  wire                _zz_181;
  wire                _zz_182;
  wire                _zz_183;
  wire                _zz_184;
  wire                _zz_185;
  wire                _zz_186;
  wire                _zz_187;
  wire                _zz_188;
  wire                _zz_189;
  wire                _zz_190;
  wire                _zz_191;
  wire                _zz_192;
  wire                _zz_193;
  wire                _zz_194;
  wire                _zz_195;
  wire                _zz_196;
  wire                _zz_197;
  wire                _zz_198;
  wire                _zz_199;
  wire                _zz_200;
  wire                _zz_201;
  wire                _zz_202;
  wire                _zz_203;
  wire                _zz_204;
  wire                _zz_205;
  wire                _zz_206;
  wire                _zz_207;
  wire                _zz_208;
  wire                _zz_209;
  wire                _zz_210;
  wire                _zz_211;
  wire                _zz_212;
  wire                _zz_213;
  wire                _zz_214;
  wire                _zz_215;
  wire                _zz_216;
  wire                _zz_217;
  wire                _zz_218;
  wire                _zz_219;
  wire                _zz_220;
  wire                _zz_221;
  wire                _zz_222;
  wire                _zz_223;
  wire                _zz_224;
  wire                _zz_225;
  wire                _zz_226;
  wire                _zz_227;
  wire                _zz_228;
  wire                _zz_229;
  wire                _zz_230;
  wire                _zz_231;
  wire                _zz_232;
  wire                _zz_233;
  wire                _zz_234;
  wire                _zz_235;
  wire                _zz_236;
  wire                _zz_237;
  wire                _zz_238;
  wire                _zz_239;
  wire                _zz_240;
  wire                _zz_241;
  wire                _zz_242;
  wire                _zz_243;
  wire                _zz_244;
  wire                _zz_245;
  wire                _zz_246;
  wire                _zz_247;
  wire                _zz_248;
  wire                _zz_249;
  wire                _zz_250;
  wire                _zz_251;
  wire                _zz_252;
  wire                _zz_253;
  wire                _zz_254;
  wire                _zz_255;
  wire                _zz_256;
  wire                _zz_257;
  wire                _zz_258;
  wire                when_DCache_l217;
  wire                when_DCache_l224;
  wire                when_DCache_l227;
  wire                when_DCache_l232;
  wire                when_DCache_l237;
  wire                when_DCache_l240;
  wire                _zz_cache_hit_1;
  wire                _zz_cache_mru_1;
  wire       [127:0]  _zz_259;
  wire                _zz_260;
  wire                _zz_261;
  wire                _zz_262;
  wire                _zz_263;
  wire                _zz_264;
  wire                _zz_265;
  wire                _zz_266;
  wire                _zz_267;
  wire                _zz_268;
  wire                _zz_269;
  wire                _zz_270;
  wire                _zz_271;
  wire                _zz_272;
  wire                _zz_273;
  wire                _zz_274;
  wire                _zz_275;
  wire                _zz_276;
  wire                _zz_277;
  wire                _zz_278;
  wire                _zz_279;
  wire                _zz_280;
  wire                _zz_281;
  wire                _zz_282;
  wire                _zz_283;
  wire                _zz_284;
  wire                _zz_285;
  wire                _zz_286;
  wire                _zz_287;
  wire                _zz_288;
  wire                _zz_289;
  wire                _zz_290;
  wire                _zz_291;
  wire                _zz_292;
  wire                _zz_293;
  wire                _zz_294;
  wire                _zz_295;
  wire                _zz_296;
  wire                _zz_297;
  wire                _zz_298;
  wire                _zz_299;
  wire                _zz_300;
  wire                _zz_301;
  wire                _zz_302;
  wire                _zz_303;
  wire                _zz_304;
  wire                _zz_305;
  wire                _zz_306;
  wire                _zz_307;
  wire                _zz_308;
  wire                _zz_309;
  wire                _zz_310;
  wire                _zz_311;
  wire                _zz_312;
  wire                _zz_313;
  wire                _zz_314;
  wire                _zz_315;
  wire                _zz_316;
  wire                _zz_317;
  wire                _zz_318;
  wire                _zz_319;
  wire                _zz_320;
  wire                _zz_321;
  wire                _zz_322;
  wire                _zz_323;
  wire                _zz_324;
  wire                _zz_325;
  wire                _zz_326;
  wire                _zz_327;
  wire                _zz_328;
  wire                _zz_329;
  wire                _zz_330;
  wire                _zz_331;
  wire                _zz_332;
  wire                _zz_333;
  wire                _zz_334;
  wire                _zz_335;
  wire                _zz_336;
  wire                _zz_337;
  wire                _zz_338;
  wire                _zz_339;
  wire                _zz_340;
  wire                _zz_341;
  wire                _zz_342;
  wire                _zz_343;
  wire                _zz_344;
  wire                _zz_345;
  wire                _zz_346;
  wire                _zz_347;
  wire                _zz_348;
  wire                _zz_349;
  wire                _zz_350;
  wire                _zz_351;
  wire                _zz_352;
  wire                _zz_353;
  wire                _zz_354;
  wire                _zz_355;
  wire                _zz_356;
  wire                _zz_357;
  wire                _zz_358;
  wire                _zz_359;
  wire                _zz_360;
  wire                _zz_361;
  wire                _zz_362;
  wire                _zz_363;
  wire                _zz_364;
  wire                _zz_365;
  wire                _zz_366;
  wire                _zz_367;
  wire                _zz_368;
  wire                _zz_369;
  wire                _zz_370;
  wire                _zz_371;
  wire                _zz_372;
  wire                _zz_373;
  wire                _zz_374;
  wire                _zz_375;
  wire                _zz_376;
  wire                _zz_377;
  wire                _zz_378;
  wire                _zz_379;
  wire                _zz_380;
  wire                _zz_381;
  wire                _zz_382;
  wire                _zz_383;
  wire                _zz_384;
  wire                _zz_385;
  wire                _zz_386;
  wire                _zz_387;
  wire                when_DCache_l181_1;
  reg        [7:0]    _zz_sram_1_ports_cmd_payload_wen;
  wire                when_DCache_l188_1;
  wire                when_DCache_l195_1;
  wire       [127:0]  _zz_388;
  wire                _zz_389;
  wire                _zz_390;
  wire                _zz_391;
  wire                _zz_392;
  wire                _zz_393;
  wire                _zz_394;
  wire                _zz_395;
  wire                _zz_396;
  wire                _zz_397;
  wire                _zz_398;
  wire                _zz_399;
  wire                _zz_400;
  wire                _zz_401;
  wire                _zz_402;
  wire                _zz_403;
  wire                _zz_404;
  wire                _zz_405;
  wire                _zz_406;
  wire                _zz_407;
  wire                _zz_408;
  wire                _zz_409;
  wire                _zz_410;
  wire                _zz_411;
  wire                _zz_412;
  wire                _zz_413;
  wire                _zz_414;
  wire                _zz_415;
  wire                _zz_416;
  wire                _zz_417;
  wire                _zz_418;
  wire                _zz_419;
  wire                _zz_420;
  wire                _zz_421;
  wire                _zz_422;
  wire                _zz_423;
  wire                _zz_424;
  wire                _zz_425;
  wire                _zz_426;
  wire                _zz_427;
  wire                _zz_428;
  wire                _zz_429;
  wire                _zz_430;
  wire                _zz_431;
  wire                _zz_432;
  wire                _zz_433;
  wire                _zz_434;
  wire                _zz_435;
  wire                _zz_436;
  wire                _zz_437;
  wire                _zz_438;
  wire                _zz_439;
  wire                _zz_440;
  wire                _zz_441;
  wire                _zz_442;
  wire                _zz_443;
  wire                _zz_444;
  wire                _zz_445;
  wire                _zz_446;
  wire                _zz_447;
  wire                _zz_448;
  wire                _zz_449;
  wire                _zz_450;
  wire                _zz_451;
  wire                _zz_452;
  wire                _zz_453;
  wire                _zz_454;
  wire                _zz_455;
  wire                _zz_456;
  wire                _zz_457;
  wire                _zz_458;
  wire                _zz_459;
  wire                _zz_460;
  wire                _zz_461;
  wire                _zz_462;
  wire                _zz_463;
  wire                _zz_464;
  wire                _zz_465;
  wire                _zz_466;
  wire                _zz_467;
  wire                _zz_468;
  wire                _zz_469;
  wire                _zz_470;
  wire                _zz_471;
  wire                _zz_472;
  wire                _zz_473;
  wire                _zz_474;
  wire                _zz_475;
  wire                _zz_476;
  wire                _zz_477;
  wire                _zz_478;
  wire                _zz_479;
  wire                _zz_480;
  wire                _zz_481;
  wire                _zz_482;
  wire                _zz_483;
  wire                _zz_484;
  wire                _zz_485;
  wire                _zz_486;
  wire                _zz_487;
  wire                _zz_488;
  wire                _zz_489;
  wire                _zz_490;
  wire                _zz_491;
  wire                _zz_492;
  wire                _zz_493;
  wire                _zz_494;
  wire                _zz_495;
  wire                _zz_496;
  wire                _zz_497;
  wire                _zz_498;
  wire                _zz_499;
  wire                _zz_500;
  wire                _zz_501;
  wire                _zz_502;
  wire                _zz_503;
  wire                _zz_504;
  wire                _zz_505;
  wire                _zz_506;
  wire                _zz_507;
  wire                _zz_508;
  wire                _zz_509;
  wire                _zz_510;
  wire                _zz_511;
  wire                _zz_512;
  wire                _zz_513;
  wire                _zz_514;
  wire                _zz_515;
  wire                _zz_516;
  wire                when_DCache_l217_1;
  wire                when_DCache_l224_1;
  wire                when_DCache_l227_1;
  wire                when_DCache_l232_1;
  wire                when_DCache_l237_1;
  wire                when_DCache_l240_1;
  wire                _zz_cache_hit_2;
  wire                _zz_cache_mru_2;
  wire       [127:0]  _zz_517;
  wire                _zz_518;
  wire                _zz_519;
  wire                _zz_520;
  wire                _zz_521;
  wire                _zz_522;
  wire                _zz_523;
  wire                _zz_524;
  wire                _zz_525;
  wire                _zz_526;
  wire                _zz_527;
  wire                _zz_528;
  wire                _zz_529;
  wire                _zz_530;
  wire                _zz_531;
  wire                _zz_532;
  wire                _zz_533;
  wire                _zz_534;
  wire                _zz_535;
  wire                _zz_536;
  wire                _zz_537;
  wire                _zz_538;
  wire                _zz_539;
  wire                _zz_540;
  wire                _zz_541;
  wire                _zz_542;
  wire                _zz_543;
  wire                _zz_544;
  wire                _zz_545;
  wire                _zz_546;
  wire                _zz_547;
  wire                _zz_548;
  wire                _zz_549;
  wire                _zz_550;
  wire                _zz_551;
  wire                _zz_552;
  wire                _zz_553;
  wire                _zz_554;
  wire                _zz_555;
  wire                _zz_556;
  wire                _zz_557;
  wire                _zz_558;
  wire                _zz_559;
  wire                _zz_560;
  wire                _zz_561;
  wire                _zz_562;
  wire                _zz_563;
  wire                _zz_564;
  wire                _zz_565;
  wire                _zz_566;
  wire                _zz_567;
  wire                _zz_568;
  wire                _zz_569;
  wire                _zz_570;
  wire                _zz_571;
  wire                _zz_572;
  wire                _zz_573;
  wire                _zz_574;
  wire                _zz_575;
  wire                _zz_576;
  wire                _zz_577;
  wire                _zz_578;
  wire                _zz_579;
  wire                _zz_580;
  wire                _zz_581;
  wire                _zz_582;
  wire                _zz_583;
  wire                _zz_584;
  wire                _zz_585;
  wire                _zz_586;
  wire                _zz_587;
  wire                _zz_588;
  wire                _zz_589;
  wire                _zz_590;
  wire                _zz_591;
  wire                _zz_592;
  wire                _zz_593;
  wire                _zz_594;
  wire                _zz_595;
  wire                _zz_596;
  wire                _zz_597;
  wire                _zz_598;
  wire                _zz_599;
  wire                _zz_600;
  wire                _zz_601;
  wire                _zz_602;
  wire                _zz_603;
  wire                _zz_604;
  wire                _zz_605;
  wire                _zz_606;
  wire                _zz_607;
  wire                _zz_608;
  wire                _zz_609;
  wire                _zz_610;
  wire                _zz_611;
  wire                _zz_612;
  wire                _zz_613;
  wire                _zz_614;
  wire                _zz_615;
  wire                _zz_616;
  wire                _zz_617;
  wire                _zz_618;
  wire                _zz_619;
  wire                _zz_620;
  wire                _zz_621;
  wire                _zz_622;
  wire                _zz_623;
  wire                _zz_624;
  wire                _zz_625;
  wire                _zz_626;
  wire                _zz_627;
  wire                _zz_628;
  wire                _zz_629;
  wire                _zz_630;
  wire                _zz_631;
  wire                _zz_632;
  wire                _zz_633;
  wire                _zz_634;
  wire                _zz_635;
  wire                _zz_636;
  wire                _zz_637;
  wire                _zz_638;
  wire                _zz_639;
  wire                _zz_640;
  wire                _zz_641;
  wire                _zz_642;
  wire                _zz_643;
  wire                _zz_644;
  wire                _zz_645;
  wire                when_DCache_l181_2;
  reg        [7:0]    _zz_sram_2_ports_cmd_payload_wen;
  wire                when_DCache_l188_2;
  wire                when_DCache_l195_2;
  wire       [127:0]  _zz_646;
  wire                _zz_647;
  wire                _zz_648;
  wire                _zz_649;
  wire                _zz_650;
  wire                _zz_651;
  wire                _zz_652;
  wire                _zz_653;
  wire                _zz_654;
  wire                _zz_655;
  wire                _zz_656;
  wire                _zz_657;
  wire                _zz_658;
  wire                _zz_659;
  wire                _zz_660;
  wire                _zz_661;
  wire                _zz_662;
  wire                _zz_663;
  wire                _zz_664;
  wire                _zz_665;
  wire                _zz_666;
  wire                _zz_667;
  wire                _zz_668;
  wire                _zz_669;
  wire                _zz_670;
  wire                _zz_671;
  wire                _zz_672;
  wire                _zz_673;
  wire                _zz_674;
  wire                _zz_675;
  wire                _zz_676;
  wire                _zz_677;
  wire                _zz_678;
  wire                _zz_679;
  wire                _zz_680;
  wire                _zz_681;
  wire                _zz_682;
  wire                _zz_683;
  wire                _zz_684;
  wire                _zz_685;
  wire                _zz_686;
  wire                _zz_687;
  wire                _zz_688;
  wire                _zz_689;
  wire                _zz_690;
  wire                _zz_691;
  wire                _zz_692;
  wire                _zz_693;
  wire                _zz_694;
  wire                _zz_695;
  wire                _zz_696;
  wire                _zz_697;
  wire                _zz_698;
  wire                _zz_699;
  wire                _zz_700;
  wire                _zz_701;
  wire                _zz_702;
  wire                _zz_703;
  wire                _zz_704;
  wire                _zz_705;
  wire                _zz_706;
  wire                _zz_707;
  wire                _zz_708;
  wire                _zz_709;
  wire                _zz_710;
  wire                _zz_711;
  wire                _zz_712;
  wire                _zz_713;
  wire                _zz_714;
  wire                _zz_715;
  wire                _zz_716;
  wire                _zz_717;
  wire                _zz_718;
  wire                _zz_719;
  wire                _zz_720;
  wire                _zz_721;
  wire                _zz_722;
  wire                _zz_723;
  wire                _zz_724;
  wire                _zz_725;
  wire                _zz_726;
  wire                _zz_727;
  wire                _zz_728;
  wire                _zz_729;
  wire                _zz_730;
  wire                _zz_731;
  wire                _zz_732;
  wire                _zz_733;
  wire                _zz_734;
  wire                _zz_735;
  wire                _zz_736;
  wire                _zz_737;
  wire                _zz_738;
  wire                _zz_739;
  wire                _zz_740;
  wire                _zz_741;
  wire                _zz_742;
  wire                _zz_743;
  wire                _zz_744;
  wire                _zz_745;
  wire                _zz_746;
  wire                _zz_747;
  wire                _zz_748;
  wire                _zz_749;
  wire                _zz_750;
  wire                _zz_751;
  wire                _zz_752;
  wire                _zz_753;
  wire                _zz_754;
  wire                _zz_755;
  wire                _zz_756;
  wire                _zz_757;
  wire                _zz_758;
  wire                _zz_759;
  wire                _zz_760;
  wire                _zz_761;
  wire                _zz_762;
  wire                _zz_763;
  wire                _zz_764;
  wire                _zz_765;
  wire                _zz_766;
  wire                _zz_767;
  wire                _zz_768;
  wire                _zz_769;
  wire                _zz_770;
  wire                _zz_771;
  wire                _zz_772;
  wire                _zz_773;
  wire                _zz_774;
  wire                when_DCache_l217_2;
  wire                when_DCache_l224_2;
  wire                when_DCache_l227_2;
  wire                when_DCache_l232_2;
  wire                when_DCache_l237_2;
  wire                when_DCache_l240_2;
  wire                _zz_cache_hit_3;
  wire                _zz_cache_mru_3;
  wire       [127:0]  _zz_775;
  wire                _zz_776;
  wire                _zz_777;
  wire                _zz_778;
  wire                _zz_779;
  wire                _zz_780;
  wire                _zz_781;
  wire                _zz_782;
  wire                _zz_783;
  wire                _zz_784;
  wire                _zz_785;
  wire                _zz_786;
  wire                _zz_787;
  wire                _zz_788;
  wire                _zz_789;
  wire                _zz_790;
  wire                _zz_791;
  wire                _zz_792;
  wire                _zz_793;
  wire                _zz_794;
  wire                _zz_795;
  wire                _zz_796;
  wire                _zz_797;
  wire                _zz_798;
  wire                _zz_799;
  wire                _zz_800;
  wire                _zz_801;
  wire                _zz_802;
  wire                _zz_803;
  wire                _zz_804;
  wire                _zz_805;
  wire                _zz_806;
  wire                _zz_807;
  wire                _zz_808;
  wire                _zz_809;
  wire                _zz_810;
  wire                _zz_811;
  wire                _zz_812;
  wire                _zz_813;
  wire                _zz_814;
  wire                _zz_815;
  wire                _zz_816;
  wire                _zz_817;
  wire                _zz_818;
  wire                _zz_819;
  wire                _zz_820;
  wire                _zz_821;
  wire                _zz_822;
  wire                _zz_823;
  wire                _zz_824;
  wire                _zz_825;
  wire                _zz_826;
  wire                _zz_827;
  wire                _zz_828;
  wire                _zz_829;
  wire                _zz_830;
  wire                _zz_831;
  wire                _zz_832;
  wire                _zz_833;
  wire                _zz_834;
  wire                _zz_835;
  wire                _zz_836;
  wire                _zz_837;
  wire                _zz_838;
  wire                _zz_839;
  wire                _zz_840;
  wire                _zz_841;
  wire                _zz_842;
  wire                _zz_843;
  wire                _zz_844;
  wire                _zz_845;
  wire                _zz_846;
  wire                _zz_847;
  wire                _zz_848;
  wire                _zz_849;
  wire                _zz_850;
  wire                _zz_851;
  wire                _zz_852;
  wire                _zz_853;
  wire                _zz_854;
  wire                _zz_855;
  wire                _zz_856;
  wire                _zz_857;
  wire                _zz_858;
  wire                _zz_859;
  wire                _zz_860;
  wire                _zz_861;
  wire                _zz_862;
  wire                _zz_863;
  wire                _zz_864;
  wire                _zz_865;
  wire                _zz_866;
  wire                _zz_867;
  wire                _zz_868;
  wire                _zz_869;
  wire                _zz_870;
  wire                _zz_871;
  wire                _zz_872;
  wire                _zz_873;
  wire                _zz_874;
  wire                _zz_875;
  wire                _zz_876;
  wire                _zz_877;
  wire                _zz_878;
  wire                _zz_879;
  wire                _zz_880;
  wire                _zz_881;
  wire                _zz_882;
  wire                _zz_883;
  wire                _zz_884;
  wire                _zz_885;
  wire                _zz_886;
  wire                _zz_887;
  wire                _zz_888;
  wire                _zz_889;
  wire                _zz_890;
  wire                _zz_891;
  wire                _zz_892;
  wire                _zz_893;
  wire                _zz_894;
  wire                _zz_895;
  wire                _zz_896;
  wire                _zz_897;
  wire                _zz_898;
  wire                _zz_899;
  wire                _zz_900;
  wire                _zz_901;
  wire                _zz_902;
  wire                _zz_903;
  wire                when_DCache_l181_3;
  reg        [7:0]    _zz_sram_3_ports_cmd_payload_wen;
  wire                when_DCache_l188_3;
  wire                when_DCache_l195_3;
  wire       [127:0]  _zz_904;
  wire                _zz_905;
  wire                _zz_906;
  wire                _zz_907;
  wire                _zz_908;
  wire                _zz_909;
  wire                _zz_910;
  wire                _zz_911;
  wire                _zz_912;
  wire                _zz_913;
  wire                _zz_914;
  wire                _zz_915;
  wire                _zz_916;
  wire                _zz_917;
  wire                _zz_918;
  wire                _zz_919;
  wire                _zz_920;
  wire                _zz_921;
  wire                _zz_922;
  wire                _zz_923;
  wire                _zz_924;
  wire                _zz_925;
  wire                _zz_926;
  wire                _zz_927;
  wire                _zz_928;
  wire                _zz_929;
  wire                _zz_930;
  wire                _zz_931;
  wire                _zz_932;
  wire                _zz_933;
  wire                _zz_934;
  wire                _zz_935;
  wire                _zz_936;
  wire                _zz_937;
  wire                _zz_938;
  wire                _zz_939;
  wire                _zz_940;
  wire                _zz_941;
  wire                _zz_942;
  wire                _zz_943;
  wire                _zz_944;
  wire                _zz_945;
  wire                _zz_946;
  wire                _zz_947;
  wire                _zz_948;
  wire                _zz_949;
  wire                _zz_950;
  wire                _zz_951;
  wire                _zz_952;
  wire                _zz_953;
  wire                _zz_954;
  wire                _zz_955;
  wire                _zz_956;
  wire                _zz_957;
  wire                _zz_958;
  wire                _zz_959;
  wire                _zz_960;
  wire                _zz_961;
  wire                _zz_962;
  wire                _zz_963;
  wire                _zz_964;
  wire                _zz_965;
  wire                _zz_966;
  wire                _zz_967;
  wire                _zz_968;
  wire                _zz_969;
  wire                _zz_970;
  wire                _zz_971;
  wire                _zz_972;
  wire                _zz_973;
  wire                _zz_974;
  wire                _zz_975;
  wire                _zz_976;
  wire                _zz_977;
  wire                _zz_978;
  wire                _zz_979;
  wire                _zz_980;
  wire                _zz_981;
  wire                _zz_982;
  wire                _zz_983;
  wire                _zz_984;
  wire                _zz_985;
  wire                _zz_986;
  wire                _zz_987;
  wire                _zz_988;
  wire                _zz_989;
  wire                _zz_990;
  wire                _zz_991;
  wire                _zz_992;
  wire                _zz_993;
  wire                _zz_994;
  wire                _zz_995;
  wire                _zz_996;
  wire                _zz_997;
  wire                _zz_998;
  wire                _zz_999;
  wire                _zz_1000;
  wire                _zz_1001;
  wire                _zz_1002;
  wire                _zz_1003;
  wire                _zz_1004;
  wire                _zz_1005;
  wire                _zz_1006;
  wire                _zz_1007;
  wire                _zz_1008;
  wire                _zz_1009;
  wire                _zz_1010;
  wire                _zz_1011;
  wire                _zz_1012;
  wire                _zz_1013;
  wire                _zz_1014;
  wire                _zz_1015;
  wire                _zz_1016;
  wire                _zz_1017;
  wire                _zz_1018;
  wire                _zz_1019;
  wire                _zz_1020;
  wire                _zz_1021;
  wire                _zz_1022;
  wire                _zz_1023;
  wire                _zz_1024;
  wire                _zz_1025;
  wire                _zz_1026;
  wire                _zz_1027;
  wire                _zz_1028;
  wire                _zz_1029;
  wire                _zz_1030;
  wire                _zz_1031;
  wire                _zz_1032;
  wire                when_DCache_l217_3;
  wire                when_DCache_l224_3;
  wire                when_DCache_l227_3;
  wire                when_DCache_l232_3;
  wire                when_DCache_l237_3;
  wire                when_DCache_l240_3;
  wire       [511:0]  _zz_cpu_rsp_payload_data;
  wire       [511:0]  _zz_cpu_rsp_payload_data_1;
  function [7:0] zz__zz_sram_0_ports_cmd_payload_wen(input dummy);
    begin
      zz__zz_sram_0_ports_cmd_payload_wen = 8'h0;
      zz__zz_sram_0_ports_cmd_payload_wen[0] = 1'b1;
    end
  endfunction
  wire [7:0] _zz_1033;
  function [7:0] zz__zz_sram_1_ports_cmd_payload_wen(input dummy);
    begin
      zz__zz_sram_1_ports_cmd_payload_wen = 8'h0;
      zz__zz_sram_1_ports_cmd_payload_wen[0] = 1'b1;
    end
  endfunction
  wire [7:0] _zz_1034;
  function [7:0] zz__zz_sram_2_ports_cmd_payload_wen(input dummy);
    begin
      zz__zz_sram_2_ports_cmd_payload_wen = 8'h0;
      zz__zz_sram_2_ports_cmd_payload_wen[0] = 1'b1;
    end
  endfunction
  wire [7:0] _zz_1035;
  function [7:0] zz__zz_sram_3_ports_cmd_payload_wen(input dummy);
    begin
      zz__zz_sram_3_ports_cmd_payload_wen = 8'h0;
      zz__zz_sram_3_ports_cmd_payload_wen[0] = 1'b1;
    end
  endfunction
  wire [7:0] _zz_1036;

  assign _zz_flush_cnt_valueNext_1 = flush_cnt_willIncrement;
  assign _zz_flush_cnt_valueNext = {6'd0, _zz_flush_cnt_valueNext_1};
  assign _zz_next_level_data_cnt_valueNext_1 = next_level_data_cnt_willIncrement;
  assign _zz_next_level_data_cnt_valueNext = {2'd0, _zz_next_level_data_cnt_valueNext_1};
  assign _zz_next_level_wstrb = (7'h0 / 4'b1000);
  assign _zz__zz_cache_hit_gnt_0_3 = (_zz_cache_hit_gnt_0_2 - _zz__zz_cache_hit_gnt_0_3_1);
  assign _zz__zz_cache_hit_gnt_0_3_2 = {_zz_cache_hit_gnt_0[3],{_zz_cache_hit_gnt_0[2],{_zz_cache_hit_gnt_0[1],_zz_cache_hit_gnt_0[0]}}};
  assign _zz__zz_cache_hit_gnt_0_3_1 = {4'd0, _zz__zz_cache_hit_gnt_0_3_2};
  assign _zz__zz_cache_invld_gnt_0_3 = (_zz_cache_invld_gnt_0_2 - _zz__zz_cache_invld_gnt_0_3_1);
  assign _zz__zz_cache_invld_gnt_0_3_2 = {_zz_cache_invld_gnt_0[3],{_zz_cache_invld_gnt_0[2],{_zz_cache_invld_gnt_0[1],_zz_cache_invld_gnt_0[0]}}};
  assign _zz__zz_cache_invld_gnt_0_3_1 = {4'd0, _zz__zz_cache_invld_gnt_0_3_2};
  assign _zz__zz_cache_victim_gnt_0_3 = (_zz_cache_victim_gnt_0_2 - _zz__zz_cache_victim_gnt_0_3_1);
  assign _zz__zz_cache_victim_gnt_0_3_2 = {_zz_cache_victim_gnt_0[3],{_zz_cache_victim_gnt_0[2],{_zz_cache_victim_gnt_0[1],_zz_cache_victim_gnt_0[0]}}};
  assign _zz__zz_cache_victim_gnt_0_3_1 = {4'd0, _zz__zz_cache_victim_gnt_0_3_2};
  assign _zz_sram_0_ports_cmd_payload_wdata = (cpu_bank_index * 7'h40);
  assign _zz_sram_0_ports_cmd_payload_wstrb = (_zz_sram_0_ports_cmd_payload_wstrb_1 / 4'b1000);
  assign _zz_sram_0_ports_cmd_payload_wstrb_1 = (cpu_bank_index * 7'h40);
  assign _zz_sram_0_ports_cmd_payload_wen_1 = (next_level_data_cnt_value * 1'b1);
  assign _zz_sram_0_ports_cmd_payload_wdata_1 = (next_level_data_cnt_value * 7'h40);
  assign _zz_sram_0_ports_cmd_payload_wstrb_2 = (_zz_sram_0_ports_cmd_payload_wstrb_3 / 4'b1000);
  assign _zz_sram_0_ports_cmd_payload_wstrb_3 = (next_level_data_cnt_value * 7'h40);
  assign _zz_sram_1_ports_cmd_payload_wdata = (cpu_bank_index * 7'h40);
  assign _zz_sram_1_ports_cmd_payload_wstrb = (_zz_sram_1_ports_cmd_payload_wstrb_1 / 4'b1000);
  assign _zz_sram_1_ports_cmd_payload_wstrb_1 = (cpu_bank_index * 7'h40);
  assign _zz_sram_1_ports_cmd_payload_wen_1 = (next_level_data_cnt_value * 1'b1);
  assign _zz_sram_1_ports_cmd_payload_wdata_1 = (next_level_data_cnt_value * 7'h40);
  assign _zz_sram_1_ports_cmd_payload_wstrb_2 = (_zz_sram_1_ports_cmd_payload_wstrb_3 / 4'b1000);
  assign _zz_sram_1_ports_cmd_payload_wstrb_3 = (next_level_data_cnt_value * 7'h40);
  assign _zz_sram_2_ports_cmd_payload_wdata = (cpu_bank_index * 7'h40);
  assign _zz_sram_2_ports_cmd_payload_wstrb = (_zz_sram_2_ports_cmd_payload_wstrb_1 / 4'b1000);
  assign _zz_sram_2_ports_cmd_payload_wstrb_1 = (cpu_bank_index * 7'h40);
  assign _zz_sram_2_ports_cmd_payload_wen_1 = (next_level_data_cnt_value * 1'b1);
  assign _zz_sram_2_ports_cmd_payload_wdata_1 = (next_level_data_cnt_value * 7'h40);
  assign _zz_sram_2_ports_cmd_payload_wstrb_2 = (_zz_sram_2_ports_cmd_payload_wstrb_3 / 4'b1000);
  assign _zz_sram_2_ports_cmd_payload_wstrb_3 = (next_level_data_cnt_value * 7'h40);
  assign _zz_sram_3_ports_cmd_payload_wdata = (cpu_bank_index * 7'h40);
  assign _zz_sram_3_ports_cmd_payload_wstrb = (_zz_sram_3_ports_cmd_payload_wstrb_1 / 4'b1000);
  assign _zz_sram_3_ports_cmd_payload_wstrb_1 = (cpu_bank_index * 7'h40);
  assign _zz_sram_3_ports_cmd_payload_wen_1 = (next_level_data_cnt_value * 1'b1);
  assign _zz_sram_3_ports_cmd_payload_wdata_1 = (next_level_data_cnt_value * 7'h40);
  assign _zz_sram_3_ports_cmd_payload_wstrb_2 = (_zz_sram_3_ports_cmd_payload_wstrb_3 / 4'b1000);
  assign _zz_sram_3_ports_cmd_payload_wstrb_3 = (next_level_data_cnt_value * 7'h40);
  always @(*) begin
    case(cpu_set)
      7'b0000000 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_0_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_0_mru;
        _zz_cache_tag_0 = ways_0_metas_0_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_0_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_0_mru;
        _zz_cache_tag_1 = ways_1_metas_0_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_0_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_0_mru;
        _zz_cache_tag_2 = ways_2_metas_0_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_0_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_0_mru;
        _zz_cache_tag_3 = ways_3_metas_0_tag;
      end
      7'b0000001 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_1_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_1_mru;
        _zz_cache_tag_0 = ways_0_metas_1_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_1_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_1_mru;
        _zz_cache_tag_1 = ways_1_metas_1_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_1_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_1_mru;
        _zz_cache_tag_2 = ways_2_metas_1_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_1_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_1_mru;
        _zz_cache_tag_3 = ways_3_metas_1_tag;
      end
      7'b0000010 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_2_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_2_mru;
        _zz_cache_tag_0 = ways_0_metas_2_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_2_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_2_mru;
        _zz_cache_tag_1 = ways_1_metas_2_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_2_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_2_mru;
        _zz_cache_tag_2 = ways_2_metas_2_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_2_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_2_mru;
        _zz_cache_tag_3 = ways_3_metas_2_tag;
      end
      7'b0000011 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_3_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_3_mru;
        _zz_cache_tag_0 = ways_0_metas_3_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_3_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_3_mru;
        _zz_cache_tag_1 = ways_1_metas_3_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_3_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_3_mru;
        _zz_cache_tag_2 = ways_2_metas_3_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_3_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_3_mru;
        _zz_cache_tag_3 = ways_3_metas_3_tag;
      end
      7'b0000100 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_4_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_4_mru;
        _zz_cache_tag_0 = ways_0_metas_4_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_4_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_4_mru;
        _zz_cache_tag_1 = ways_1_metas_4_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_4_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_4_mru;
        _zz_cache_tag_2 = ways_2_metas_4_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_4_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_4_mru;
        _zz_cache_tag_3 = ways_3_metas_4_tag;
      end
      7'b0000101 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_5_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_5_mru;
        _zz_cache_tag_0 = ways_0_metas_5_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_5_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_5_mru;
        _zz_cache_tag_1 = ways_1_metas_5_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_5_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_5_mru;
        _zz_cache_tag_2 = ways_2_metas_5_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_5_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_5_mru;
        _zz_cache_tag_3 = ways_3_metas_5_tag;
      end
      7'b0000110 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_6_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_6_mru;
        _zz_cache_tag_0 = ways_0_metas_6_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_6_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_6_mru;
        _zz_cache_tag_1 = ways_1_metas_6_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_6_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_6_mru;
        _zz_cache_tag_2 = ways_2_metas_6_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_6_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_6_mru;
        _zz_cache_tag_3 = ways_3_metas_6_tag;
      end
      7'b0000111 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_7_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_7_mru;
        _zz_cache_tag_0 = ways_0_metas_7_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_7_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_7_mru;
        _zz_cache_tag_1 = ways_1_metas_7_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_7_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_7_mru;
        _zz_cache_tag_2 = ways_2_metas_7_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_7_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_7_mru;
        _zz_cache_tag_3 = ways_3_metas_7_tag;
      end
      7'b0001000 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_8_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_8_mru;
        _zz_cache_tag_0 = ways_0_metas_8_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_8_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_8_mru;
        _zz_cache_tag_1 = ways_1_metas_8_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_8_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_8_mru;
        _zz_cache_tag_2 = ways_2_metas_8_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_8_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_8_mru;
        _zz_cache_tag_3 = ways_3_metas_8_tag;
      end
      7'b0001001 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_9_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_9_mru;
        _zz_cache_tag_0 = ways_0_metas_9_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_9_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_9_mru;
        _zz_cache_tag_1 = ways_1_metas_9_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_9_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_9_mru;
        _zz_cache_tag_2 = ways_2_metas_9_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_9_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_9_mru;
        _zz_cache_tag_3 = ways_3_metas_9_tag;
      end
      7'b0001010 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_10_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_10_mru;
        _zz_cache_tag_0 = ways_0_metas_10_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_10_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_10_mru;
        _zz_cache_tag_1 = ways_1_metas_10_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_10_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_10_mru;
        _zz_cache_tag_2 = ways_2_metas_10_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_10_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_10_mru;
        _zz_cache_tag_3 = ways_3_metas_10_tag;
      end
      7'b0001011 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_11_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_11_mru;
        _zz_cache_tag_0 = ways_0_metas_11_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_11_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_11_mru;
        _zz_cache_tag_1 = ways_1_metas_11_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_11_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_11_mru;
        _zz_cache_tag_2 = ways_2_metas_11_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_11_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_11_mru;
        _zz_cache_tag_3 = ways_3_metas_11_tag;
      end
      7'b0001100 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_12_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_12_mru;
        _zz_cache_tag_0 = ways_0_metas_12_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_12_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_12_mru;
        _zz_cache_tag_1 = ways_1_metas_12_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_12_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_12_mru;
        _zz_cache_tag_2 = ways_2_metas_12_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_12_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_12_mru;
        _zz_cache_tag_3 = ways_3_metas_12_tag;
      end
      7'b0001101 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_13_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_13_mru;
        _zz_cache_tag_0 = ways_0_metas_13_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_13_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_13_mru;
        _zz_cache_tag_1 = ways_1_metas_13_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_13_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_13_mru;
        _zz_cache_tag_2 = ways_2_metas_13_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_13_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_13_mru;
        _zz_cache_tag_3 = ways_3_metas_13_tag;
      end
      7'b0001110 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_14_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_14_mru;
        _zz_cache_tag_0 = ways_0_metas_14_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_14_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_14_mru;
        _zz_cache_tag_1 = ways_1_metas_14_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_14_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_14_mru;
        _zz_cache_tag_2 = ways_2_metas_14_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_14_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_14_mru;
        _zz_cache_tag_3 = ways_3_metas_14_tag;
      end
      7'b0001111 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_15_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_15_mru;
        _zz_cache_tag_0 = ways_0_metas_15_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_15_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_15_mru;
        _zz_cache_tag_1 = ways_1_metas_15_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_15_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_15_mru;
        _zz_cache_tag_2 = ways_2_metas_15_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_15_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_15_mru;
        _zz_cache_tag_3 = ways_3_metas_15_tag;
      end
      7'b0010000 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_16_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_16_mru;
        _zz_cache_tag_0 = ways_0_metas_16_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_16_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_16_mru;
        _zz_cache_tag_1 = ways_1_metas_16_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_16_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_16_mru;
        _zz_cache_tag_2 = ways_2_metas_16_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_16_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_16_mru;
        _zz_cache_tag_3 = ways_3_metas_16_tag;
      end
      7'b0010001 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_17_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_17_mru;
        _zz_cache_tag_0 = ways_0_metas_17_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_17_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_17_mru;
        _zz_cache_tag_1 = ways_1_metas_17_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_17_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_17_mru;
        _zz_cache_tag_2 = ways_2_metas_17_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_17_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_17_mru;
        _zz_cache_tag_3 = ways_3_metas_17_tag;
      end
      7'b0010010 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_18_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_18_mru;
        _zz_cache_tag_0 = ways_0_metas_18_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_18_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_18_mru;
        _zz_cache_tag_1 = ways_1_metas_18_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_18_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_18_mru;
        _zz_cache_tag_2 = ways_2_metas_18_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_18_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_18_mru;
        _zz_cache_tag_3 = ways_3_metas_18_tag;
      end
      7'b0010011 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_19_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_19_mru;
        _zz_cache_tag_0 = ways_0_metas_19_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_19_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_19_mru;
        _zz_cache_tag_1 = ways_1_metas_19_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_19_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_19_mru;
        _zz_cache_tag_2 = ways_2_metas_19_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_19_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_19_mru;
        _zz_cache_tag_3 = ways_3_metas_19_tag;
      end
      7'b0010100 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_20_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_20_mru;
        _zz_cache_tag_0 = ways_0_metas_20_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_20_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_20_mru;
        _zz_cache_tag_1 = ways_1_metas_20_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_20_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_20_mru;
        _zz_cache_tag_2 = ways_2_metas_20_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_20_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_20_mru;
        _zz_cache_tag_3 = ways_3_metas_20_tag;
      end
      7'b0010101 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_21_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_21_mru;
        _zz_cache_tag_0 = ways_0_metas_21_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_21_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_21_mru;
        _zz_cache_tag_1 = ways_1_metas_21_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_21_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_21_mru;
        _zz_cache_tag_2 = ways_2_metas_21_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_21_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_21_mru;
        _zz_cache_tag_3 = ways_3_metas_21_tag;
      end
      7'b0010110 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_22_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_22_mru;
        _zz_cache_tag_0 = ways_0_metas_22_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_22_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_22_mru;
        _zz_cache_tag_1 = ways_1_metas_22_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_22_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_22_mru;
        _zz_cache_tag_2 = ways_2_metas_22_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_22_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_22_mru;
        _zz_cache_tag_3 = ways_3_metas_22_tag;
      end
      7'b0010111 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_23_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_23_mru;
        _zz_cache_tag_0 = ways_0_metas_23_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_23_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_23_mru;
        _zz_cache_tag_1 = ways_1_metas_23_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_23_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_23_mru;
        _zz_cache_tag_2 = ways_2_metas_23_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_23_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_23_mru;
        _zz_cache_tag_3 = ways_3_metas_23_tag;
      end
      7'b0011000 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_24_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_24_mru;
        _zz_cache_tag_0 = ways_0_metas_24_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_24_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_24_mru;
        _zz_cache_tag_1 = ways_1_metas_24_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_24_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_24_mru;
        _zz_cache_tag_2 = ways_2_metas_24_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_24_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_24_mru;
        _zz_cache_tag_3 = ways_3_metas_24_tag;
      end
      7'b0011001 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_25_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_25_mru;
        _zz_cache_tag_0 = ways_0_metas_25_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_25_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_25_mru;
        _zz_cache_tag_1 = ways_1_metas_25_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_25_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_25_mru;
        _zz_cache_tag_2 = ways_2_metas_25_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_25_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_25_mru;
        _zz_cache_tag_3 = ways_3_metas_25_tag;
      end
      7'b0011010 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_26_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_26_mru;
        _zz_cache_tag_0 = ways_0_metas_26_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_26_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_26_mru;
        _zz_cache_tag_1 = ways_1_metas_26_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_26_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_26_mru;
        _zz_cache_tag_2 = ways_2_metas_26_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_26_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_26_mru;
        _zz_cache_tag_3 = ways_3_metas_26_tag;
      end
      7'b0011011 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_27_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_27_mru;
        _zz_cache_tag_0 = ways_0_metas_27_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_27_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_27_mru;
        _zz_cache_tag_1 = ways_1_metas_27_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_27_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_27_mru;
        _zz_cache_tag_2 = ways_2_metas_27_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_27_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_27_mru;
        _zz_cache_tag_3 = ways_3_metas_27_tag;
      end
      7'b0011100 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_28_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_28_mru;
        _zz_cache_tag_0 = ways_0_metas_28_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_28_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_28_mru;
        _zz_cache_tag_1 = ways_1_metas_28_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_28_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_28_mru;
        _zz_cache_tag_2 = ways_2_metas_28_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_28_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_28_mru;
        _zz_cache_tag_3 = ways_3_metas_28_tag;
      end
      7'b0011101 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_29_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_29_mru;
        _zz_cache_tag_0 = ways_0_metas_29_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_29_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_29_mru;
        _zz_cache_tag_1 = ways_1_metas_29_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_29_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_29_mru;
        _zz_cache_tag_2 = ways_2_metas_29_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_29_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_29_mru;
        _zz_cache_tag_3 = ways_3_metas_29_tag;
      end
      7'b0011110 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_30_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_30_mru;
        _zz_cache_tag_0 = ways_0_metas_30_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_30_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_30_mru;
        _zz_cache_tag_1 = ways_1_metas_30_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_30_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_30_mru;
        _zz_cache_tag_2 = ways_2_metas_30_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_30_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_30_mru;
        _zz_cache_tag_3 = ways_3_metas_30_tag;
      end
      7'b0011111 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_31_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_31_mru;
        _zz_cache_tag_0 = ways_0_metas_31_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_31_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_31_mru;
        _zz_cache_tag_1 = ways_1_metas_31_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_31_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_31_mru;
        _zz_cache_tag_2 = ways_2_metas_31_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_31_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_31_mru;
        _zz_cache_tag_3 = ways_3_metas_31_tag;
      end
      7'b0100000 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_32_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_32_mru;
        _zz_cache_tag_0 = ways_0_metas_32_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_32_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_32_mru;
        _zz_cache_tag_1 = ways_1_metas_32_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_32_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_32_mru;
        _zz_cache_tag_2 = ways_2_metas_32_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_32_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_32_mru;
        _zz_cache_tag_3 = ways_3_metas_32_tag;
      end
      7'b0100001 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_33_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_33_mru;
        _zz_cache_tag_0 = ways_0_metas_33_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_33_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_33_mru;
        _zz_cache_tag_1 = ways_1_metas_33_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_33_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_33_mru;
        _zz_cache_tag_2 = ways_2_metas_33_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_33_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_33_mru;
        _zz_cache_tag_3 = ways_3_metas_33_tag;
      end
      7'b0100010 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_34_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_34_mru;
        _zz_cache_tag_0 = ways_0_metas_34_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_34_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_34_mru;
        _zz_cache_tag_1 = ways_1_metas_34_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_34_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_34_mru;
        _zz_cache_tag_2 = ways_2_metas_34_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_34_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_34_mru;
        _zz_cache_tag_3 = ways_3_metas_34_tag;
      end
      7'b0100011 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_35_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_35_mru;
        _zz_cache_tag_0 = ways_0_metas_35_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_35_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_35_mru;
        _zz_cache_tag_1 = ways_1_metas_35_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_35_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_35_mru;
        _zz_cache_tag_2 = ways_2_metas_35_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_35_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_35_mru;
        _zz_cache_tag_3 = ways_3_metas_35_tag;
      end
      7'b0100100 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_36_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_36_mru;
        _zz_cache_tag_0 = ways_0_metas_36_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_36_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_36_mru;
        _zz_cache_tag_1 = ways_1_metas_36_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_36_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_36_mru;
        _zz_cache_tag_2 = ways_2_metas_36_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_36_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_36_mru;
        _zz_cache_tag_3 = ways_3_metas_36_tag;
      end
      7'b0100101 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_37_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_37_mru;
        _zz_cache_tag_0 = ways_0_metas_37_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_37_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_37_mru;
        _zz_cache_tag_1 = ways_1_metas_37_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_37_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_37_mru;
        _zz_cache_tag_2 = ways_2_metas_37_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_37_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_37_mru;
        _zz_cache_tag_3 = ways_3_metas_37_tag;
      end
      7'b0100110 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_38_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_38_mru;
        _zz_cache_tag_0 = ways_0_metas_38_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_38_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_38_mru;
        _zz_cache_tag_1 = ways_1_metas_38_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_38_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_38_mru;
        _zz_cache_tag_2 = ways_2_metas_38_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_38_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_38_mru;
        _zz_cache_tag_3 = ways_3_metas_38_tag;
      end
      7'b0100111 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_39_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_39_mru;
        _zz_cache_tag_0 = ways_0_metas_39_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_39_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_39_mru;
        _zz_cache_tag_1 = ways_1_metas_39_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_39_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_39_mru;
        _zz_cache_tag_2 = ways_2_metas_39_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_39_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_39_mru;
        _zz_cache_tag_3 = ways_3_metas_39_tag;
      end
      7'b0101000 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_40_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_40_mru;
        _zz_cache_tag_0 = ways_0_metas_40_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_40_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_40_mru;
        _zz_cache_tag_1 = ways_1_metas_40_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_40_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_40_mru;
        _zz_cache_tag_2 = ways_2_metas_40_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_40_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_40_mru;
        _zz_cache_tag_3 = ways_3_metas_40_tag;
      end
      7'b0101001 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_41_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_41_mru;
        _zz_cache_tag_0 = ways_0_metas_41_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_41_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_41_mru;
        _zz_cache_tag_1 = ways_1_metas_41_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_41_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_41_mru;
        _zz_cache_tag_2 = ways_2_metas_41_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_41_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_41_mru;
        _zz_cache_tag_3 = ways_3_metas_41_tag;
      end
      7'b0101010 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_42_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_42_mru;
        _zz_cache_tag_0 = ways_0_metas_42_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_42_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_42_mru;
        _zz_cache_tag_1 = ways_1_metas_42_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_42_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_42_mru;
        _zz_cache_tag_2 = ways_2_metas_42_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_42_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_42_mru;
        _zz_cache_tag_3 = ways_3_metas_42_tag;
      end
      7'b0101011 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_43_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_43_mru;
        _zz_cache_tag_0 = ways_0_metas_43_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_43_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_43_mru;
        _zz_cache_tag_1 = ways_1_metas_43_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_43_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_43_mru;
        _zz_cache_tag_2 = ways_2_metas_43_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_43_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_43_mru;
        _zz_cache_tag_3 = ways_3_metas_43_tag;
      end
      7'b0101100 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_44_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_44_mru;
        _zz_cache_tag_0 = ways_0_metas_44_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_44_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_44_mru;
        _zz_cache_tag_1 = ways_1_metas_44_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_44_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_44_mru;
        _zz_cache_tag_2 = ways_2_metas_44_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_44_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_44_mru;
        _zz_cache_tag_3 = ways_3_metas_44_tag;
      end
      7'b0101101 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_45_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_45_mru;
        _zz_cache_tag_0 = ways_0_metas_45_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_45_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_45_mru;
        _zz_cache_tag_1 = ways_1_metas_45_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_45_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_45_mru;
        _zz_cache_tag_2 = ways_2_metas_45_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_45_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_45_mru;
        _zz_cache_tag_3 = ways_3_metas_45_tag;
      end
      7'b0101110 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_46_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_46_mru;
        _zz_cache_tag_0 = ways_0_metas_46_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_46_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_46_mru;
        _zz_cache_tag_1 = ways_1_metas_46_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_46_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_46_mru;
        _zz_cache_tag_2 = ways_2_metas_46_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_46_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_46_mru;
        _zz_cache_tag_3 = ways_3_metas_46_tag;
      end
      7'b0101111 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_47_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_47_mru;
        _zz_cache_tag_0 = ways_0_metas_47_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_47_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_47_mru;
        _zz_cache_tag_1 = ways_1_metas_47_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_47_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_47_mru;
        _zz_cache_tag_2 = ways_2_metas_47_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_47_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_47_mru;
        _zz_cache_tag_3 = ways_3_metas_47_tag;
      end
      7'b0110000 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_48_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_48_mru;
        _zz_cache_tag_0 = ways_0_metas_48_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_48_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_48_mru;
        _zz_cache_tag_1 = ways_1_metas_48_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_48_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_48_mru;
        _zz_cache_tag_2 = ways_2_metas_48_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_48_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_48_mru;
        _zz_cache_tag_3 = ways_3_metas_48_tag;
      end
      7'b0110001 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_49_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_49_mru;
        _zz_cache_tag_0 = ways_0_metas_49_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_49_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_49_mru;
        _zz_cache_tag_1 = ways_1_metas_49_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_49_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_49_mru;
        _zz_cache_tag_2 = ways_2_metas_49_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_49_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_49_mru;
        _zz_cache_tag_3 = ways_3_metas_49_tag;
      end
      7'b0110010 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_50_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_50_mru;
        _zz_cache_tag_0 = ways_0_metas_50_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_50_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_50_mru;
        _zz_cache_tag_1 = ways_1_metas_50_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_50_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_50_mru;
        _zz_cache_tag_2 = ways_2_metas_50_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_50_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_50_mru;
        _zz_cache_tag_3 = ways_3_metas_50_tag;
      end
      7'b0110011 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_51_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_51_mru;
        _zz_cache_tag_0 = ways_0_metas_51_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_51_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_51_mru;
        _zz_cache_tag_1 = ways_1_metas_51_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_51_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_51_mru;
        _zz_cache_tag_2 = ways_2_metas_51_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_51_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_51_mru;
        _zz_cache_tag_3 = ways_3_metas_51_tag;
      end
      7'b0110100 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_52_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_52_mru;
        _zz_cache_tag_0 = ways_0_metas_52_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_52_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_52_mru;
        _zz_cache_tag_1 = ways_1_metas_52_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_52_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_52_mru;
        _zz_cache_tag_2 = ways_2_metas_52_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_52_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_52_mru;
        _zz_cache_tag_3 = ways_3_metas_52_tag;
      end
      7'b0110101 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_53_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_53_mru;
        _zz_cache_tag_0 = ways_0_metas_53_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_53_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_53_mru;
        _zz_cache_tag_1 = ways_1_metas_53_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_53_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_53_mru;
        _zz_cache_tag_2 = ways_2_metas_53_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_53_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_53_mru;
        _zz_cache_tag_3 = ways_3_metas_53_tag;
      end
      7'b0110110 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_54_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_54_mru;
        _zz_cache_tag_0 = ways_0_metas_54_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_54_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_54_mru;
        _zz_cache_tag_1 = ways_1_metas_54_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_54_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_54_mru;
        _zz_cache_tag_2 = ways_2_metas_54_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_54_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_54_mru;
        _zz_cache_tag_3 = ways_3_metas_54_tag;
      end
      7'b0110111 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_55_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_55_mru;
        _zz_cache_tag_0 = ways_0_metas_55_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_55_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_55_mru;
        _zz_cache_tag_1 = ways_1_metas_55_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_55_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_55_mru;
        _zz_cache_tag_2 = ways_2_metas_55_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_55_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_55_mru;
        _zz_cache_tag_3 = ways_3_metas_55_tag;
      end
      7'b0111000 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_56_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_56_mru;
        _zz_cache_tag_0 = ways_0_metas_56_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_56_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_56_mru;
        _zz_cache_tag_1 = ways_1_metas_56_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_56_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_56_mru;
        _zz_cache_tag_2 = ways_2_metas_56_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_56_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_56_mru;
        _zz_cache_tag_3 = ways_3_metas_56_tag;
      end
      7'b0111001 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_57_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_57_mru;
        _zz_cache_tag_0 = ways_0_metas_57_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_57_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_57_mru;
        _zz_cache_tag_1 = ways_1_metas_57_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_57_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_57_mru;
        _zz_cache_tag_2 = ways_2_metas_57_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_57_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_57_mru;
        _zz_cache_tag_3 = ways_3_metas_57_tag;
      end
      7'b0111010 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_58_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_58_mru;
        _zz_cache_tag_0 = ways_0_metas_58_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_58_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_58_mru;
        _zz_cache_tag_1 = ways_1_metas_58_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_58_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_58_mru;
        _zz_cache_tag_2 = ways_2_metas_58_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_58_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_58_mru;
        _zz_cache_tag_3 = ways_3_metas_58_tag;
      end
      7'b0111011 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_59_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_59_mru;
        _zz_cache_tag_0 = ways_0_metas_59_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_59_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_59_mru;
        _zz_cache_tag_1 = ways_1_metas_59_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_59_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_59_mru;
        _zz_cache_tag_2 = ways_2_metas_59_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_59_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_59_mru;
        _zz_cache_tag_3 = ways_3_metas_59_tag;
      end
      7'b0111100 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_60_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_60_mru;
        _zz_cache_tag_0 = ways_0_metas_60_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_60_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_60_mru;
        _zz_cache_tag_1 = ways_1_metas_60_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_60_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_60_mru;
        _zz_cache_tag_2 = ways_2_metas_60_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_60_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_60_mru;
        _zz_cache_tag_3 = ways_3_metas_60_tag;
      end
      7'b0111101 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_61_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_61_mru;
        _zz_cache_tag_0 = ways_0_metas_61_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_61_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_61_mru;
        _zz_cache_tag_1 = ways_1_metas_61_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_61_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_61_mru;
        _zz_cache_tag_2 = ways_2_metas_61_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_61_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_61_mru;
        _zz_cache_tag_3 = ways_3_metas_61_tag;
      end
      7'b0111110 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_62_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_62_mru;
        _zz_cache_tag_0 = ways_0_metas_62_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_62_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_62_mru;
        _zz_cache_tag_1 = ways_1_metas_62_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_62_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_62_mru;
        _zz_cache_tag_2 = ways_2_metas_62_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_62_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_62_mru;
        _zz_cache_tag_3 = ways_3_metas_62_tag;
      end
      7'b0111111 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_63_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_63_mru;
        _zz_cache_tag_0 = ways_0_metas_63_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_63_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_63_mru;
        _zz_cache_tag_1 = ways_1_metas_63_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_63_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_63_mru;
        _zz_cache_tag_2 = ways_2_metas_63_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_63_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_63_mru;
        _zz_cache_tag_3 = ways_3_metas_63_tag;
      end
      7'b1000000 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_64_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_64_mru;
        _zz_cache_tag_0 = ways_0_metas_64_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_64_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_64_mru;
        _zz_cache_tag_1 = ways_1_metas_64_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_64_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_64_mru;
        _zz_cache_tag_2 = ways_2_metas_64_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_64_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_64_mru;
        _zz_cache_tag_3 = ways_3_metas_64_tag;
      end
      7'b1000001 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_65_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_65_mru;
        _zz_cache_tag_0 = ways_0_metas_65_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_65_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_65_mru;
        _zz_cache_tag_1 = ways_1_metas_65_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_65_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_65_mru;
        _zz_cache_tag_2 = ways_2_metas_65_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_65_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_65_mru;
        _zz_cache_tag_3 = ways_3_metas_65_tag;
      end
      7'b1000010 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_66_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_66_mru;
        _zz_cache_tag_0 = ways_0_metas_66_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_66_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_66_mru;
        _zz_cache_tag_1 = ways_1_metas_66_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_66_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_66_mru;
        _zz_cache_tag_2 = ways_2_metas_66_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_66_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_66_mru;
        _zz_cache_tag_3 = ways_3_metas_66_tag;
      end
      7'b1000011 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_67_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_67_mru;
        _zz_cache_tag_0 = ways_0_metas_67_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_67_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_67_mru;
        _zz_cache_tag_1 = ways_1_metas_67_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_67_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_67_mru;
        _zz_cache_tag_2 = ways_2_metas_67_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_67_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_67_mru;
        _zz_cache_tag_3 = ways_3_metas_67_tag;
      end
      7'b1000100 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_68_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_68_mru;
        _zz_cache_tag_0 = ways_0_metas_68_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_68_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_68_mru;
        _zz_cache_tag_1 = ways_1_metas_68_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_68_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_68_mru;
        _zz_cache_tag_2 = ways_2_metas_68_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_68_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_68_mru;
        _zz_cache_tag_3 = ways_3_metas_68_tag;
      end
      7'b1000101 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_69_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_69_mru;
        _zz_cache_tag_0 = ways_0_metas_69_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_69_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_69_mru;
        _zz_cache_tag_1 = ways_1_metas_69_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_69_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_69_mru;
        _zz_cache_tag_2 = ways_2_metas_69_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_69_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_69_mru;
        _zz_cache_tag_3 = ways_3_metas_69_tag;
      end
      7'b1000110 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_70_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_70_mru;
        _zz_cache_tag_0 = ways_0_metas_70_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_70_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_70_mru;
        _zz_cache_tag_1 = ways_1_metas_70_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_70_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_70_mru;
        _zz_cache_tag_2 = ways_2_metas_70_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_70_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_70_mru;
        _zz_cache_tag_3 = ways_3_metas_70_tag;
      end
      7'b1000111 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_71_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_71_mru;
        _zz_cache_tag_0 = ways_0_metas_71_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_71_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_71_mru;
        _zz_cache_tag_1 = ways_1_metas_71_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_71_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_71_mru;
        _zz_cache_tag_2 = ways_2_metas_71_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_71_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_71_mru;
        _zz_cache_tag_3 = ways_3_metas_71_tag;
      end
      7'b1001000 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_72_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_72_mru;
        _zz_cache_tag_0 = ways_0_metas_72_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_72_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_72_mru;
        _zz_cache_tag_1 = ways_1_metas_72_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_72_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_72_mru;
        _zz_cache_tag_2 = ways_2_metas_72_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_72_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_72_mru;
        _zz_cache_tag_3 = ways_3_metas_72_tag;
      end
      7'b1001001 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_73_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_73_mru;
        _zz_cache_tag_0 = ways_0_metas_73_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_73_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_73_mru;
        _zz_cache_tag_1 = ways_1_metas_73_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_73_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_73_mru;
        _zz_cache_tag_2 = ways_2_metas_73_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_73_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_73_mru;
        _zz_cache_tag_3 = ways_3_metas_73_tag;
      end
      7'b1001010 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_74_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_74_mru;
        _zz_cache_tag_0 = ways_0_metas_74_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_74_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_74_mru;
        _zz_cache_tag_1 = ways_1_metas_74_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_74_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_74_mru;
        _zz_cache_tag_2 = ways_2_metas_74_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_74_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_74_mru;
        _zz_cache_tag_3 = ways_3_metas_74_tag;
      end
      7'b1001011 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_75_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_75_mru;
        _zz_cache_tag_0 = ways_0_metas_75_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_75_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_75_mru;
        _zz_cache_tag_1 = ways_1_metas_75_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_75_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_75_mru;
        _zz_cache_tag_2 = ways_2_metas_75_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_75_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_75_mru;
        _zz_cache_tag_3 = ways_3_metas_75_tag;
      end
      7'b1001100 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_76_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_76_mru;
        _zz_cache_tag_0 = ways_0_metas_76_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_76_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_76_mru;
        _zz_cache_tag_1 = ways_1_metas_76_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_76_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_76_mru;
        _zz_cache_tag_2 = ways_2_metas_76_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_76_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_76_mru;
        _zz_cache_tag_3 = ways_3_metas_76_tag;
      end
      7'b1001101 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_77_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_77_mru;
        _zz_cache_tag_0 = ways_0_metas_77_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_77_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_77_mru;
        _zz_cache_tag_1 = ways_1_metas_77_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_77_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_77_mru;
        _zz_cache_tag_2 = ways_2_metas_77_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_77_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_77_mru;
        _zz_cache_tag_3 = ways_3_metas_77_tag;
      end
      7'b1001110 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_78_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_78_mru;
        _zz_cache_tag_0 = ways_0_metas_78_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_78_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_78_mru;
        _zz_cache_tag_1 = ways_1_metas_78_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_78_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_78_mru;
        _zz_cache_tag_2 = ways_2_metas_78_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_78_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_78_mru;
        _zz_cache_tag_3 = ways_3_metas_78_tag;
      end
      7'b1001111 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_79_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_79_mru;
        _zz_cache_tag_0 = ways_0_metas_79_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_79_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_79_mru;
        _zz_cache_tag_1 = ways_1_metas_79_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_79_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_79_mru;
        _zz_cache_tag_2 = ways_2_metas_79_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_79_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_79_mru;
        _zz_cache_tag_3 = ways_3_metas_79_tag;
      end
      7'b1010000 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_80_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_80_mru;
        _zz_cache_tag_0 = ways_0_metas_80_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_80_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_80_mru;
        _zz_cache_tag_1 = ways_1_metas_80_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_80_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_80_mru;
        _zz_cache_tag_2 = ways_2_metas_80_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_80_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_80_mru;
        _zz_cache_tag_3 = ways_3_metas_80_tag;
      end
      7'b1010001 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_81_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_81_mru;
        _zz_cache_tag_0 = ways_0_metas_81_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_81_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_81_mru;
        _zz_cache_tag_1 = ways_1_metas_81_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_81_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_81_mru;
        _zz_cache_tag_2 = ways_2_metas_81_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_81_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_81_mru;
        _zz_cache_tag_3 = ways_3_metas_81_tag;
      end
      7'b1010010 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_82_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_82_mru;
        _zz_cache_tag_0 = ways_0_metas_82_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_82_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_82_mru;
        _zz_cache_tag_1 = ways_1_metas_82_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_82_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_82_mru;
        _zz_cache_tag_2 = ways_2_metas_82_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_82_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_82_mru;
        _zz_cache_tag_3 = ways_3_metas_82_tag;
      end
      7'b1010011 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_83_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_83_mru;
        _zz_cache_tag_0 = ways_0_metas_83_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_83_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_83_mru;
        _zz_cache_tag_1 = ways_1_metas_83_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_83_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_83_mru;
        _zz_cache_tag_2 = ways_2_metas_83_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_83_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_83_mru;
        _zz_cache_tag_3 = ways_3_metas_83_tag;
      end
      7'b1010100 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_84_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_84_mru;
        _zz_cache_tag_0 = ways_0_metas_84_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_84_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_84_mru;
        _zz_cache_tag_1 = ways_1_metas_84_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_84_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_84_mru;
        _zz_cache_tag_2 = ways_2_metas_84_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_84_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_84_mru;
        _zz_cache_tag_3 = ways_3_metas_84_tag;
      end
      7'b1010101 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_85_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_85_mru;
        _zz_cache_tag_0 = ways_0_metas_85_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_85_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_85_mru;
        _zz_cache_tag_1 = ways_1_metas_85_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_85_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_85_mru;
        _zz_cache_tag_2 = ways_2_metas_85_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_85_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_85_mru;
        _zz_cache_tag_3 = ways_3_metas_85_tag;
      end
      7'b1010110 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_86_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_86_mru;
        _zz_cache_tag_0 = ways_0_metas_86_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_86_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_86_mru;
        _zz_cache_tag_1 = ways_1_metas_86_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_86_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_86_mru;
        _zz_cache_tag_2 = ways_2_metas_86_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_86_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_86_mru;
        _zz_cache_tag_3 = ways_3_metas_86_tag;
      end
      7'b1010111 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_87_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_87_mru;
        _zz_cache_tag_0 = ways_0_metas_87_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_87_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_87_mru;
        _zz_cache_tag_1 = ways_1_metas_87_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_87_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_87_mru;
        _zz_cache_tag_2 = ways_2_metas_87_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_87_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_87_mru;
        _zz_cache_tag_3 = ways_3_metas_87_tag;
      end
      7'b1011000 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_88_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_88_mru;
        _zz_cache_tag_0 = ways_0_metas_88_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_88_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_88_mru;
        _zz_cache_tag_1 = ways_1_metas_88_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_88_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_88_mru;
        _zz_cache_tag_2 = ways_2_metas_88_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_88_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_88_mru;
        _zz_cache_tag_3 = ways_3_metas_88_tag;
      end
      7'b1011001 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_89_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_89_mru;
        _zz_cache_tag_0 = ways_0_metas_89_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_89_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_89_mru;
        _zz_cache_tag_1 = ways_1_metas_89_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_89_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_89_mru;
        _zz_cache_tag_2 = ways_2_metas_89_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_89_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_89_mru;
        _zz_cache_tag_3 = ways_3_metas_89_tag;
      end
      7'b1011010 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_90_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_90_mru;
        _zz_cache_tag_0 = ways_0_metas_90_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_90_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_90_mru;
        _zz_cache_tag_1 = ways_1_metas_90_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_90_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_90_mru;
        _zz_cache_tag_2 = ways_2_metas_90_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_90_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_90_mru;
        _zz_cache_tag_3 = ways_3_metas_90_tag;
      end
      7'b1011011 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_91_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_91_mru;
        _zz_cache_tag_0 = ways_0_metas_91_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_91_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_91_mru;
        _zz_cache_tag_1 = ways_1_metas_91_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_91_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_91_mru;
        _zz_cache_tag_2 = ways_2_metas_91_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_91_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_91_mru;
        _zz_cache_tag_3 = ways_3_metas_91_tag;
      end
      7'b1011100 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_92_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_92_mru;
        _zz_cache_tag_0 = ways_0_metas_92_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_92_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_92_mru;
        _zz_cache_tag_1 = ways_1_metas_92_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_92_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_92_mru;
        _zz_cache_tag_2 = ways_2_metas_92_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_92_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_92_mru;
        _zz_cache_tag_3 = ways_3_metas_92_tag;
      end
      7'b1011101 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_93_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_93_mru;
        _zz_cache_tag_0 = ways_0_metas_93_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_93_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_93_mru;
        _zz_cache_tag_1 = ways_1_metas_93_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_93_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_93_mru;
        _zz_cache_tag_2 = ways_2_metas_93_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_93_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_93_mru;
        _zz_cache_tag_3 = ways_3_metas_93_tag;
      end
      7'b1011110 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_94_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_94_mru;
        _zz_cache_tag_0 = ways_0_metas_94_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_94_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_94_mru;
        _zz_cache_tag_1 = ways_1_metas_94_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_94_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_94_mru;
        _zz_cache_tag_2 = ways_2_metas_94_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_94_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_94_mru;
        _zz_cache_tag_3 = ways_3_metas_94_tag;
      end
      7'b1011111 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_95_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_95_mru;
        _zz_cache_tag_0 = ways_0_metas_95_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_95_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_95_mru;
        _zz_cache_tag_1 = ways_1_metas_95_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_95_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_95_mru;
        _zz_cache_tag_2 = ways_2_metas_95_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_95_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_95_mru;
        _zz_cache_tag_3 = ways_3_metas_95_tag;
      end
      7'b1100000 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_96_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_96_mru;
        _zz_cache_tag_0 = ways_0_metas_96_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_96_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_96_mru;
        _zz_cache_tag_1 = ways_1_metas_96_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_96_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_96_mru;
        _zz_cache_tag_2 = ways_2_metas_96_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_96_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_96_mru;
        _zz_cache_tag_3 = ways_3_metas_96_tag;
      end
      7'b1100001 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_97_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_97_mru;
        _zz_cache_tag_0 = ways_0_metas_97_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_97_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_97_mru;
        _zz_cache_tag_1 = ways_1_metas_97_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_97_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_97_mru;
        _zz_cache_tag_2 = ways_2_metas_97_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_97_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_97_mru;
        _zz_cache_tag_3 = ways_3_metas_97_tag;
      end
      7'b1100010 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_98_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_98_mru;
        _zz_cache_tag_0 = ways_0_metas_98_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_98_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_98_mru;
        _zz_cache_tag_1 = ways_1_metas_98_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_98_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_98_mru;
        _zz_cache_tag_2 = ways_2_metas_98_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_98_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_98_mru;
        _zz_cache_tag_3 = ways_3_metas_98_tag;
      end
      7'b1100011 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_99_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_99_mru;
        _zz_cache_tag_0 = ways_0_metas_99_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_99_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_99_mru;
        _zz_cache_tag_1 = ways_1_metas_99_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_99_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_99_mru;
        _zz_cache_tag_2 = ways_2_metas_99_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_99_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_99_mru;
        _zz_cache_tag_3 = ways_3_metas_99_tag;
      end
      7'b1100100 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_100_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_100_mru;
        _zz_cache_tag_0 = ways_0_metas_100_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_100_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_100_mru;
        _zz_cache_tag_1 = ways_1_metas_100_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_100_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_100_mru;
        _zz_cache_tag_2 = ways_2_metas_100_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_100_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_100_mru;
        _zz_cache_tag_3 = ways_3_metas_100_tag;
      end
      7'b1100101 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_101_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_101_mru;
        _zz_cache_tag_0 = ways_0_metas_101_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_101_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_101_mru;
        _zz_cache_tag_1 = ways_1_metas_101_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_101_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_101_mru;
        _zz_cache_tag_2 = ways_2_metas_101_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_101_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_101_mru;
        _zz_cache_tag_3 = ways_3_metas_101_tag;
      end
      7'b1100110 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_102_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_102_mru;
        _zz_cache_tag_0 = ways_0_metas_102_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_102_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_102_mru;
        _zz_cache_tag_1 = ways_1_metas_102_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_102_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_102_mru;
        _zz_cache_tag_2 = ways_2_metas_102_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_102_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_102_mru;
        _zz_cache_tag_3 = ways_3_metas_102_tag;
      end
      7'b1100111 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_103_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_103_mru;
        _zz_cache_tag_0 = ways_0_metas_103_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_103_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_103_mru;
        _zz_cache_tag_1 = ways_1_metas_103_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_103_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_103_mru;
        _zz_cache_tag_2 = ways_2_metas_103_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_103_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_103_mru;
        _zz_cache_tag_3 = ways_3_metas_103_tag;
      end
      7'b1101000 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_104_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_104_mru;
        _zz_cache_tag_0 = ways_0_metas_104_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_104_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_104_mru;
        _zz_cache_tag_1 = ways_1_metas_104_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_104_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_104_mru;
        _zz_cache_tag_2 = ways_2_metas_104_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_104_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_104_mru;
        _zz_cache_tag_3 = ways_3_metas_104_tag;
      end
      7'b1101001 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_105_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_105_mru;
        _zz_cache_tag_0 = ways_0_metas_105_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_105_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_105_mru;
        _zz_cache_tag_1 = ways_1_metas_105_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_105_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_105_mru;
        _zz_cache_tag_2 = ways_2_metas_105_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_105_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_105_mru;
        _zz_cache_tag_3 = ways_3_metas_105_tag;
      end
      7'b1101010 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_106_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_106_mru;
        _zz_cache_tag_0 = ways_0_metas_106_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_106_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_106_mru;
        _zz_cache_tag_1 = ways_1_metas_106_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_106_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_106_mru;
        _zz_cache_tag_2 = ways_2_metas_106_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_106_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_106_mru;
        _zz_cache_tag_3 = ways_3_metas_106_tag;
      end
      7'b1101011 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_107_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_107_mru;
        _zz_cache_tag_0 = ways_0_metas_107_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_107_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_107_mru;
        _zz_cache_tag_1 = ways_1_metas_107_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_107_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_107_mru;
        _zz_cache_tag_2 = ways_2_metas_107_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_107_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_107_mru;
        _zz_cache_tag_3 = ways_3_metas_107_tag;
      end
      7'b1101100 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_108_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_108_mru;
        _zz_cache_tag_0 = ways_0_metas_108_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_108_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_108_mru;
        _zz_cache_tag_1 = ways_1_metas_108_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_108_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_108_mru;
        _zz_cache_tag_2 = ways_2_metas_108_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_108_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_108_mru;
        _zz_cache_tag_3 = ways_3_metas_108_tag;
      end
      7'b1101101 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_109_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_109_mru;
        _zz_cache_tag_0 = ways_0_metas_109_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_109_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_109_mru;
        _zz_cache_tag_1 = ways_1_metas_109_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_109_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_109_mru;
        _zz_cache_tag_2 = ways_2_metas_109_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_109_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_109_mru;
        _zz_cache_tag_3 = ways_3_metas_109_tag;
      end
      7'b1101110 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_110_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_110_mru;
        _zz_cache_tag_0 = ways_0_metas_110_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_110_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_110_mru;
        _zz_cache_tag_1 = ways_1_metas_110_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_110_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_110_mru;
        _zz_cache_tag_2 = ways_2_metas_110_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_110_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_110_mru;
        _zz_cache_tag_3 = ways_3_metas_110_tag;
      end
      7'b1101111 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_111_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_111_mru;
        _zz_cache_tag_0 = ways_0_metas_111_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_111_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_111_mru;
        _zz_cache_tag_1 = ways_1_metas_111_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_111_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_111_mru;
        _zz_cache_tag_2 = ways_2_metas_111_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_111_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_111_mru;
        _zz_cache_tag_3 = ways_3_metas_111_tag;
      end
      7'b1110000 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_112_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_112_mru;
        _zz_cache_tag_0 = ways_0_metas_112_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_112_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_112_mru;
        _zz_cache_tag_1 = ways_1_metas_112_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_112_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_112_mru;
        _zz_cache_tag_2 = ways_2_metas_112_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_112_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_112_mru;
        _zz_cache_tag_3 = ways_3_metas_112_tag;
      end
      7'b1110001 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_113_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_113_mru;
        _zz_cache_tag_0 = ways_0_metas_113_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_113_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_113_mru;
        _zz_cache_tag_1 = ways_1_metas_113_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_113_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_113_mru;
        _zz_cache_tag_2 = ways_2_metas_113_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_113_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_113_mru;
        _zz_cache_tag_3 = ways_3_metas_113_tag;
      end
      7'b1110010 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_114_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_114_mru;
        _zz_cache_tag_0 = ways_0_metas_114_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_114_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_114_mru;
        _zz_cache_tag_1 = ways_1_metas_114_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_114_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_114_mru;
        _zz_cache_tag_2 = ways_2_metas_114_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_114_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_114_mru;
        _zz_cache_tag_3 = ways_3_metas_114_tag;
      end
      7'b1110011 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_115_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_115_mru;
        _zz_cache_tag_0 = ways_0_metas_115_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_115_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_115_mru;
        _zz_cache_tag_1 = ways_1_metas_115_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_115_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_115_mru;
        _zz_cache_tag_2 = ways_2_metas_115_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_115_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_115_mru;
        _zz_cache_tag_3 = ways_3_metas_115_tag;
      end
      7'b1110100 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_116_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_116_mru;
        _zz_cache_tag_0 = ways_0_metas_116_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_116_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_116_mru;
        _zz_cache_tag_1 = ways_1_metas_116_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_116_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_116_mru;
        _zz_cache_tag_2 = ways_2_metas_116_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_116_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_116_mru;
        _zz_cache_tag_3 = ways_3_metas_116_tag;
      end
      7'b1110101 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_117_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_117_mru;
        _zz_cache_tag_0 = ways_0_metas_117_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_117_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_117_mru;
        _zz_cache_tag_1 = ways_1_metas_117_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_117_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_117_mru;
        _zz_cache_tag_2 = ways_2_metas_117_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_117_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_117_mru;
        _zz_cache_tag_3 = ways_3_metas_117_tag;
      end
      7'b1110110 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_118_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_118_mru;
        _zz_cache_tag_0 = ways_0_metas_118_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_118_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_118_mru;
        _zz_cache_tag_1 = ways_1_metas_118_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_118_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_118_mru;
        _zz_cache_tag_2 = ways_2_metas_118_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_118_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_118_mru;
        _zz_cache_tag_3 = ways_3_metas_118_tag;
      end
      7'b1110111 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_119_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_119_mru;
        _zz_cache_tag_0 = ways_0_metas_119_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_119_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_119_mru;
        _zz_cache_tag_1 = ways_1_metas_119_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_119_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_119_mru;
        _zz_cache_tag_2 = ways_2_metas_119_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_119_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_119_mru;
        _zz_cache_tag_3 = ways_3_metas_119_tag;
      end
      7'b1111000 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_120_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_120_mru;
        _zz_cache_tag_0 = ways_0_metas_120_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_120_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_120_mru;
        _zz_cache_tag_1 = ways_1_metas_120_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_120_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_120_mru;
        _zz_cache_tag_2 = ways_2_metas_120_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_120_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_120_mru;
        _zz_cache_tag_3 = ways_3_metas_120_tag;
      end
      7'b1111001 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_121_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_121_mru;
        _zz_cache_tag_0 = ways_0_metas_121_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_121_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_121_mru;
        _zz_cache_tag_1 = ways_1_metas_121_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_121_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_121_mru;
        _zz_cache_tag_2 = ways_2_metas_121_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_121_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_121_mru;
        _zz_cache_tag_3 = ways_3_metas_121_tag;
      end
      7'b1111010 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_122_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_122_mru;
        _zz_cache_tag_0 = ways_0_metas_122_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_122_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_122_mru;
        _zz_cache_tag_1 = ways_1_metas_122_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_122_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_122_mru;
        _zz_cache_tag_2 = ways_2_metas_122_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_122_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_122_mru;
        _zz_cache_tag_3 = ways_3_metas_122_tag;
      end
      7'b1111011 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_123_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_123_mru;
        _zz_cache_tag_0 = ways_0_metas_123_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_123_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_123_mru;
        _zz_cache_tag_1 = ways_1_metas_123_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_123_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_123_mru;
        _zz_cache_tag_2 = ways_2_metas_123_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_123_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_123_mru;
        _zz_cache_tag_3 = ways_3_metas_123_tag;
      end
      7'b1111100 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_124_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_124_mru;
        _zz_cache_tag_0 = ways_0_metas_124_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_124_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_124_mru;
        _zz_cache_tag_1 = ways_1_metas_124_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_124_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_124_mru;
        _zz_cache_tag_2 = ways_2_metas_124_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_124_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_124_mru;
        _zz_cache_tag_3 = ways_3_metas_124_tag;
      end
      7'b1111101 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_125_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_125_mru;
        _zz_cache_tag_0 = ways_0_metas_125_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_125_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_125_mru;
        _zz_cache_tag_1 = ways_1_metas_125_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_125_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_125_mru;
        _zz_cache_tag_2 = ways_2_metas_125_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_125_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_125_mru;
        _zz_cache_tag_3 = ways_3_metas_125_tag;
      end
      7'b1111110 : begin
        _zz__zz_cache_hit_0 = ways_0_metas_126_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_126_mru;
        _zz_cache_tag_0 = ways_0_metas_126_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_126_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_126_mru;
        _zz_cache_tag_1 = ways_1_metas_126_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_126_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_126_mru;
        _zz_cache_tag_2 = ways_2_metas_126_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_126_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_126_mru;
        _zz_cache_tag_3 = ways_3_metas_126_tag;
      end
      default : begin
        _zz__zz_cache_hit_0 = ways_0_metas_127_vld;
        _zz__zz_cache_mru_0 = ways_0_metas_127_mru;
        _zz_cache_tag_0 = ways_0_metas_127_tag;
        _zz__zz_cache_hit_1 = ways_1_metas_127_vld;
        _zz__zz_cache_mru_1 = ways_1_metas_127_mru;
        _zz_cache_tag_1 = ways_1_metas_127_tag;
        _zz__zz_cache_hit_2 = ways_2_metas_127_vld;
        _zz__zz_cache_mru_2 = ways_2_metas_127_mru;
        _zz_cache_tag_2 = ways_2_metas_127_tag;
        _zz__zz_cache_hit_3 = ways_3_metas_127_vld;
        _zz__zz_cache_mru_3 = ways_3_metas_127_mru;
        _zz_cache_tag_3 = ways_3_metas_127_tag;
      end
    endcase
  end

  always @(*) begin
    case(hit_id)
      2'b00 : begin
        _zz__zz_cpu_rsp_payload_data = sram_banks_data_0;
        _zz_cpu_rsp_valid = sram_banks_valid_0;
      end
      2'b01 : begin
        _zz__zz_cpu_rsp_payload_data = sram_banks_data_1;
        _zz_cpu_rsp_valid = sram_banks_valid_1;
      end
      2'b10 : begin
        _zz__zz_cpu_rsp_payload_data = sram_banks_data_2;
        _zz_cpu_rsp_valid = sram_banks_valid_2;
      end
      default : begin
        _zz__zz_cpu_rsp_payload_data = sram_banks_data_3;
        _zz_cpu_rsp_valid = sram_banks_valid_3;
      end
    endcase
  end

  always @(*) begin
    case(evict_id_miss)
      2'b00 : begin
        _zz__zz_cpu_rsp_payload_data_1 = sram_banks_data_0;
        _zz_cpu_rsp_valid_1 = sram_banks_valid_0;
      end
      2'b01 : begin
        _zz__zz_cpu_rsp_payload_data_1 = sram_banks_data_1;
        _zz_cpu_rsp_valid_1 = sram_banks_valid_1;
      end
      2'b10 : begin
        _zz__zz_cpu_rsp_payload_data_1 = sram_banks_data_2;
        _zz_cpu_rsp_valid_1 = sram_banks_valid_2;
      end
      default : begin
        _zz__zz_cpu_rsp_payload_data_1 = sram_banks_data_3;
        _zz_cpu_rsp_valid_1 = sram_banks_valid_3;
      end
    endcase
  end

  always @(*) begin
    case(cpu_bank_index)
      3'b000 : begin
        _zz_cpu_rsp_payload_data_2 = _zz_cpu_rsp_payload_data[63 : 0];
        _zz_cpu_rsp_payload_data_3 = _zz_cpu_rsp_payload_data_1[63 : 0];
      end
      3'b001 : begin
        _zz_cpu_rsp_payload_data_2 = _zz_cpu_rsp_payload_data[127 : 64];
        _zz_cpu_rsp_payload_data_3 = _zz_cpu_rsp_payload_data_1[127 : 64];
      end
      3'b010 : begin
        _zz_cpu_rsp_payload_data_2 = _zz_cpu_rsp_payload_data[191 : 128];
        _zz_cpu_rsp_payload_data_3 = _zz_cpu_rsp_payload_data_1[191 : 128];
      end
      3'b011 : begin
        _zz_cpu_rsp_payload_data_2 = _zz_cpu_rsp_payload_data[255 : 192];
        _zz_cpu_rsp_payload_data_3 = _zz_cpu_rsp_payload_data_1[255 : 192];
      end
      3'b100 : begin
        _zz_cpu_rsp_payload_data_2 = _zz_cpu_rsp_payload_data[319 : 256];
        _zz_cpu_rsp_payload_data_3 = _zz_cpu_rsp_payload_data_1[319 : 256];
      end
      3'b101 : begin
        _zz_cpu_rsp_payload_data_2 = _zz_cpu_rsp_payload_data[383 : 320];
        _zz_cpu_rsp_payload_data_3 = _zz_cpu_rsp_payload_data_1[383 : 320];
      end
      3'b110 : begin
        _zz_cpu_rsp_payload_data_2 = _zz_cpu_rsp_payload_data[447 : 384];
        _zz_cpu_rsp_payload_data_3 = _zz_cpu_rsp_payload_data_1[447 : 384];
      end
      default : begin
        _zz_cpu_rsp_payload_data_2 = _zz_cpu_rsp_payload_data[511 : 448];
        _zz_cpu_rsp_payload_data_3 = _zz_cpu_rsp_payload_data_1[511 : 448];
      end
    endcase
  end

  assign mru_full = (&{cache_mru_3,{cache_mru_2,{cache_mru_1,cache_mru_0}}});
  assign cpu_cmd_fire = (cpu_cmd_valid && cpu_cmd_ready);
  assign is_hit = ((|{cache_hit_3,{cache_hit_2,{cache_hit_1,cache_hit_0}}}) && cpu_cmd_fire);
  assign cpu_cmd_fire_1 = (cpu_cmd_valid && cpu_cmd_ready);
  assign is_miss = ((! (|{cache_hit_3,{cache_hit_2,{cache_hit_1,cache_hit_0}}})) && cpu_cmd_fire_1);
  assign is_diff = (! (|{cache_victim_3,{cache_victim_2,{cache_victim_1,cache_victim_0}}}));
  assign cpu_cmd_fire_2 = (cpu_cmd_valid && cpu_cmd_ready);
  assign is_write = (cpu_cmd_fire_2 && cpu_cmd_payload_wen);
  always @(*) begin
    flush_cnt_willIncrement = 1'b0;
    if(!when_DCache_l149) begin
      if(flush_busy) begin
        flush_cnt_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    flush_cnt_willClear = 1'b0;
    if(when_DCache_l149) begin
      flush_cnt_willClear = 1'b1;
    end
  end

  assign flush_cnt_willOverflowIfInc = (flush_cnt_value == 7'h7f);
  assign flush_cnt_willOverflow = (flush_cnt_willOverflowIfInc && flush_cnt_willIncrement);
  always @(*) begin
    flush_cnt_valueNext = (flush_cnt_value + _zz_flush_cnt_valueNext);
    if(flush_cnt_willClear) begin
      flush_cnt_valueNext = 7'h0;
    end
  end

  assign flush_done = (flush_busy && (flush_cnt_value == 7'h7f));
  assign cpu_tag = cpu_cmd_payload_addr[63 : 13];
  assign cpu_set = cpu_cmd_payload_addr[12 : 6];
  assign cpu_bank_addr = cpu_cmd_payload_addr[12 : 6];
  assign cpu_bank_index = cpu_cmd_payload_addr[5 : 3];
  always @(*) begin
    next_level_data_cnt_willIncrement = 1'b0;
    if(!when_DCache_l131) begin
      if(!next_level_rdone) begin
        if(next_level_rvalid) begin
          next_level_data_cnt_willIncrement = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    next_level_data_cnt_willClear = 1'b0;
    if(when_DCache_l131) begin
      next_level_data_cnt_willClear = 1'b1;
    end else begin
      if(next_level_rdone) begin
        next_level_data_cnt_willClear = 1'b1;
      end
    end
  end

  assign next_level_data_cnt_willOverflowIfInc = (next_level_data_cnt_value == 3'b111);
  assign next_level_data_cnt_willOverflow = (next_level_data_cnt_willOverflowIfInc && next_level_data_cnt_willIncrement);
  always @(*) begin
    next_level_data_cnt_valueNext = (next_level_data_cnt_value + _zz_next_level_data_cnt_valueNext);
    if(next_level_data_cnt_willClear) begin
      next_level_data_cnt_valueNext = 3'b000;
    end
  end

  assign next_level_bank_addr = cpu_cmd_payload_addr[12 : 6];
  assign next_level_rvalid = (next_level_rsp_valid && next_level_rsp_payload_rvalid);
  assign next_level_wstrb_tmp = cpu_cmd_payload_wstrb;
  assign next_level_wdata_tmp = cpu_cmd_payload_wdata;
  assign next_level_wstrb = (next_level_wstrb_tmp <<< _zz_next_level_wstrb);
  assign next_level_wdata = (next_level_wdata_tmp <<< 7'h0);
  assign when_DCache_l123 = (is_miss || is_write);
  assign when_DCache_l131 = (is_miss && (! is_write));
  assign when_DCache_l149 = (flush_busy && (flush_cnt_value == 7'h7f));
  assign _zz_cache_hit_gnt_0 = 4'b0001;
  assign _zz_cache_hit_gnt_0_1 = {cache_hit_3,{cache_hit_2,{cache_hit_1,cache_hit_0}}};
  assign _zz_cache_hit_gnt_0_2 = {_zz_cache_hit_gnt_0_1,_zz_cache_hit_gnt_0_1};
  assign _zz_cache_hit_gnt_0_3 = (_zz_cache_hit_gnt_0_2 & (~ _zz__zz_cache_hit_gnt_0_3));
  assign _zz_cache_hit_gnt_0_4 = (_zz_cache_hit_gnt_0_3[7 : 4] | _zz_cache_hit_gnt_0_3[3 : 0]);
  assign cache_hit_gnt_0 = _zz_cache_hit_gnt_0_4[0];
  assign cache_hit_gnt_1 = _zz_cache_hit_gnt_0_4[1];
  assign cache_hit_gnt_2 = _zz_cache_hit_gnt_0_4[2];
  assign cache_hit_gnt_3 = _zz_cache_hit_gnt_0_4[3];
  assign _zz_cache_invld_gnt_0 = 4'b0001;
  assign _zz_cache_invld_gnt_0_1 = {cache_invld_3,{cache_invld_2,{cache_invld_1,cache_invld_0}}};
  assign _zz_cache_invld_gnt_0_2 = {_zz_cache_invld_gnt_0_1,_zz_cache_invld_gnt_0_1};
  assign _zz_cache_invld_gnt_0_3 = (_zz_cache_invld_gnt_0_2 & (~ _zz__zz_cache_invld_gnt_0_3));
  assign _zz_cache_invld_gnt_0_4 = (_zz_cache_invld_gnt_0_3[7 : 4] | _zz_cache_invld_gnt_0_3[3 : 0]);
  assign cache_invld_gnt_0 = _zz_cache_invld_gnt_0_4[0];
  assign cache_invld_gnt_1 = _zz_cache_invld_gnt_0_4[1];
  assign cache_invld_gnt_2 = _zz_cache_invld_gnt_0_4[2];
  assign cache_invld_gnt_3 = _zz_cache_invld_gnt_0_4[3];
  assign _zz_cache_victim_gnt_0 = 4'b0001;
  assign _zz_cache_victim_gnt_0_1 = {cache_victim_3,{cache_victim_2,{cache_victim_1,cache_victim_0}}};
  assign _zz_cache_victim_gnt_0_2 = {_zz_cache_victim_gnt_0_1,_zz_cache_victim_gnt_0_1};
  assign _zz_cache_victim_gnt_0_3 = (_zz_cache_victim_gnt_0_2 & (~ _zz__zz_cache_victim_gnt_0_3));
  assign _zz_cache_victim_gnt_0_4 = (_zz_cache_victim_gnt_0_3[7 : 4] | _zz_cache_victim_gnt_0_3[3 : 0]);
  assign cache_victim_gnt_0 = _zz_cache_victim_gnt_0_4[0];
  assign cache_victim_gnt_1 = _zz_cache_victim_gnt_0_4[1];
  assign cache_victim_gnt_2 = _zz_cache_victim_gnt_0_4[2];
  assign cache_victim_gnt_3 = _zz_cache_victim_gnt_0_4[3];
  assign _zz_hit_id = (cache_hit_gnt_1 || cache_hit_gnt_3);
  assign _zz_hit_id_1 = (cache_hit_gnt_2 || cache_hit_gnt_3);
  assign hit_id = {_zz_hit_id_1,_zz_hit_id};
  assign _zz_invld_id = (cache_invld_gnt_1 || cache_invld_gnt_3);
  assign _zz_invld_id_1 = (cache_invld_gnt_2 || cache_invld_gnt_3);
  assign invld_id = {_zz_invld_id_1,_zz_invld_id};
  assign _zz_victim_id = (cache_victim_gnt_1 || cache_victim_gnt_3);
  assign _zz_victim_id_1 = (cache_victim_gnt_2 || cache_victim_gnt_3);
  assign victim_id = {_zz_victim_id_1,_zz_victim_id};
  assign evict_id = (is_diff ? invld_id : victim_id);
  assign _zz_cache_hit_0 = _zz__zz_cache_hit_0;
  assign _zz_cache_mru_0 = _zz__zz_cache_mru_0;
  assign _zz_1 = ({127'd0,1'b1} <<< cpu_set);
  assign _zz_2 = _zz_1[0];
  assign _zz_3 = _zz_1[1];
  assign _zz_4 = _zz_1[2];
  assign _zz_5 = _zz_1[3];
  assign _zz_6 = _zz_1[4];
  assign _zz_7 = _zz_1[5];
  assign _zz_8 = _zz_1[6];
  assign _zz_9 = _zz_1[7];
  assign _zz_10 = _zz_1[8];
  assign _zz_11 = _zz_1[9];
  assign _zz_12 = _zz_1[10];
  assign _zz_13 = _zz_1[11];
  assign _zz_14 = _zz_1[12];
  assign _zz_15 = _zz_1[13];
  assign _zz_16 = _zz_1[14];
  assign _zz_17 = _zz_1[15];
  assign _zz_18 = _zz_1[16];
  assign _zz_19 = _zz_1[17];
  assign _zz_20 = _zz_1[18];
  assign _zz_21 = _zz_1[19];
  assign _zz_22 = _zz_1[20];
  assign _zz_23 = _zz_1[21];
  assign _zz_24 = _zz_1[22];
  assign _zz_25 = _zz_1[23];
  assign _zz_26 = _zz_1[24];
  assign _zz_27 = _zz_1[25];
  assign _zz_28 = _zz_1[26];
  assign _zz_29 = _zz_1[27];
  assign _zz_30 = _zz_1[28];
  assign _zz_31 = _zz_1[29];
  assign _zz_32 = _zz_1[30];
  assign _zz_33 = _zz_1[31];
  assign _zz_34 = _zz_1[32];
  assign _zz_35 = _zz_1[33];
  assign _zz_36 = _zz_1[34];
  assign _zz_37 = _zz_1[35];
  assign _zz_38 = _zz_1[36];
  assign _zz_39 = _zz_1[37];
  assign _zz_40 = _zz_1[38];
  assign _zz_41 = _zz_1[39];
  assign _zz_42 = _zz_1[40];
  assign _zz_43 = _zz_1[41];
  assign _zz_44 = _zz_1[42];
  assign _zz_45 = _zz_1[43];
  assign _zz_46 = _zz_1[44];
  assign _zz_47 = _zz_1[45];
  assign _zz_48 = _zz_1[46];
  assign _zz_49 = _zz_1[47];
  assign _zz_50 = _zz_1[48];
  assign _zz_51 = _zz_1[49];
  assign _zz_52 = _zz_1[50];
  assign _zz_53 = _zz_1[51];
  assign _zz_54 = _zz_1[52];
  assign _zz_55 = _zz_1[53];
  assign _zz_56 = _zz_1[54];
  assign _zz_57 = _zz_1[55];
  assign _zz_58 = _zz_1[56];
  assign _zz_59 = _zz_1[57];
  assign _zz_60 = _zz_1[58];
  assign _zz_61 = _zz_1[59];
  assign _zz_62 = _zz_1[60];
  assign _zz_63 = _zz_1[61];
  assign _zz_64 = _zz_1[62];
  assign _zz_65 = _zz_1[63];
  assign _zz_66 = _zz_1[64];
  assign _zz_67 = _zz_1[65];
  assign _zz_68 = _zz_1[66];
  assign _zz_69 = _zz_1[67];
  assign _zz_70 = _zz_1[68];
  assign _zz_71 = _zz_1[69];
  assign _zz_72 = _zz_1[70];
  assign _zz_73 = _zz_1[71];
  assign _zz_74 = _zz_1[72];
  assign _zz_75 = _zz_1[73];
  assign _zz_76 = _zz_1[74];
  assign _zz_77 = _zz_1[75];
  assign _zz_78 = _zz_1[76];
  assign _zz_79 = _zz_1[77];
  assign _zz_80 = _zz_1[78];
  assign _zz_81 = _zz_1[79];
  assign _zz_82 = _zz_1[80];
  assign _zz_83 = _zz_1[81];
  assign _zz_84 = _zz_1[82];
  assign _zz_85 = _zz_1[83];
  assign _zz_86 = _zz_1[84];
  assign _zz_87 = _zz_1[85];
  assign _zz_88 = _zz_1[86];
  assign _zz_89 = _zz_1[87];
  assign _zz_90 = _zz_1[88];
  assign _zz_91 = _zz_1[89];
  assign _zz_92 = _zz_1[90];
  assign _zz_93 = _zz_1[91];
  assign _zz_94 = _zz_1[92];
  assign _zz_95 = _zz_1[93];
  assign _zz_96 = _zz_1[94];
  assign _zz_97 = _zz_1[95];
  assign _zz_98 = _zz_1[96];
  assign _zz_99 = _zz_1[97];
  assign _zz_100 = _zz_1[98];
  assign _zz_101 = _zz_1[99];
  assign _zz_102 = _zz_1[100];
  assign _zz_103 = _zz_1[101];
  assign _zz_104 = _zz_1[102];
  assign _zz_105 = _zz_1[103];
  assign _zz_106 = _zz_1[104];
  assign _zz_107 = _zz_1[105];
  assign _zz_108 = _zz_1[106];
  assign _zz_109 = _zz_1[107];
  assign _zz_110 = _zz_1[108];
  assign _zz_111 = _zz_1[109];
  assign _zz_112 = _zz_1[110];
  assign _zz_113 = _zz_1[111];
  assign _zz_114 = _zz_1[112];
  assign _zz_115 = _zz_1[113];
  assign _zz_116 = _zz_1[114];
  assign _zz_117 = _zz_1[115];
  assign _zz_118 = _zz_1[116];
  assign _zz_119 = _zz_1[117];
  assign _zz_120 = _zz_1[118];
  assign _zz_121 = _zz_1[119];
  assign _zz_122 = _zz_1[120];
  assign _zz_123 = _zz_1[121];
  assign _zz_124 = _zz_1[122];
  assign _zz_125 = _zz_1[123];
  assign _zz_126 = _zz_1[124];
  assign _zz_127 = _zz_1[125];
  assign _zz_128 = _zz_1[126];
  assign _zz_129 = _zz_1[127];
  assign cache_tag_0 = _zz_cache_tag_0;
  assign cache_hit_0 = ((cache_tag_0 == cpu_tag) && _zz_cache_hit_0);
  assign cache_mru_0 = _zz_cache_mru_0;
  assign cache_invld_0 = (! _zz_cache_hit_0);
  assign cache_lru_0 = (! _zz_cache_mru_0);
  assign cache_victim_0 = (cache_invld_0 && cache_lru_0);
  assign sram_banks_data_0 = sram_0_ports_rsp_payload_data;
  assign sram_banks_valid_0 = sram_0_ports_rsp_valid;
  assign when_DCache_l181 = (is_hit && (2'b00 == hit_id));
  always @(*) begin
    if(when_DCache_l181) begin
      sram_0_ports_cmd_payload_addr = cpu_bank_addr;
    end else begin
      if(when_DCache_l188) begin
        sram_0_ports_cmd_payload_addr = cpu_bank_addr;
      end else begin
        if(when_DCache_l195) begin
          sram_0_ports_cmd_payload_addr = next_level_bank_addr;
        end else begin
          sram_0_ports_cmd_payload_addr = 7'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l181) begin
      sram_0_ports_cmd_valid = 1'b1;
    end else begin
      if(when_DCache_l188) begin
        sram_0_ports_cmd_valid = 1'b1;
      end else begin
        if(when_DCache_l195) begin
          sram_0_ports_cmd_valid = 1'b1;
        end else begin
          sram_0_ports_cmd_valid = 1'b0;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l181) begin
      sram_0_ports_cmd_payload_wen = ({7'h0,cpu_cmd_payload_wen} <<< cpu_bank_index);
    end else begin
      if(when_DCache_l188) begin
        sram_0_ports_cmd_payload_wen = 8'h0;
      end else begin
        if(when_DCache_l195) begin
          sram_0_ports_cmd_payload_wen = (_zz_sram_0_ports_cmd_payload_wen <<< _zz_sram_0_ports_cmd_payload_wen_1);
        end else begin
          sram_0_ports_cmd_payload_wen = 8'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l181) begin
      sram_0_ports_cmd_payload_wdata = ({448'h0,cpu_cmd_payload_wdata} <<< _zz_sram_0_ports_cmd_payload_wdata);
    end else begin
      if(when_DCache_l188) begin
        sram_0_ports_cmd_payload_wdata = 512'h0;
      end else begin
        if(when_DCache_l195) begin
          sram_0_ports_cmd_payload_wdata = ({448'h0,next_level_rsp_payload_data} <<< _zz_sram_0_ports_cmd_payload_wdata_1);
        end else begin
          sram_0_ports_cmd_payload_wdata = 512'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l181) begin
      sram_0_ports_cmd_payload_wstrb = ({56'h0,cpu_cmd_payload_wstrb} <<< _zz_sram_0_ports_cmd_payload_wstrb);
    end else begin
      if(when_DCache_l188) begin
        sram_0_ports_cmd_payload_wstrb = 64'h0;
      end else begin
        if(when_DCache_l195) begin
          sram_0_ports_cmd_payload_wstrb = ({56'h0,8'hff} <<< _zz_sram_0_ports_cmd_payload_wstrb_2);
        end else begin
          sram_0_ports_cmd_payload_wstrb = 64'h0;
        end
      end
    end
  end

  assign _zz_1033 = zz__zz_sram_0_ports_cmd_payload_wen(1'b0);
  always @(*) _zz_sram_0_ports_cmd_payload_wen = _zz_1033;
  assign when_DCache_l188 = ((next_level_rdone && (! is_write)) && (2'b00 == evict_id_miss));
  assign when_DCache_l195 = (next_level_rvalid && (2'b00 == evict_id_miss));
  assign _zz_130 = ({127'd0,1'b1} <<< flush_cnt_value);
  assign _zz_131 = _zz_130[0];
  assign _zz_132 = _zz_130[1];
  assign _zz_133 = _zz_130[2];
  assign _zz_134 = _zz_130[3];
  assign _zz_135 = _zz_130[4];
  assign _zz_136 = _zz_130[5];
  assign _zz_137 = _zz_130[6];
  assign _zz_138 = _zz_130[7];
  assign _zz_139 = _zz_130[8];
  assign _zz_140 = _zz_130[9];
  assign _zz_141 = _zz_130[10];
  assign _zz_142 = _zz_130[11];
  assign _zz_143 = _zz_130[12];
  assign _zz_144 = _zz_130[13];
  assign _zz_145 = _zz_130[14];
  assign _zz_146 = _zz_130[15];
  assign _zz_147 = _zz_130[16];
  assign _zz_148 = _zz_130[17];
  assign _zz_149 = _zz_130[18];
  assign _zz_150 = _zz_130[19];
  assign _zz_151 = _zz_130[20];
  assign _zz_152 = _zz_130[21];
  assign _zz_153 = _zz_130[22];
  assign _zz_154 = _zz_130[23];
  assign _zz_155 = _zz_130[24];
  assign _zz_156 = _zz_130[25];
  assign _zz_157 = _zz_130[26];
  assign _zz_158 = _zz_130[27];
  assign _zz_159 = _zz_130[28];
  assign _zz_160 = _zz_130[29];
  assign _zz_161 = _zz_130[30];
  assign _zz_162 = _zz_130[31];
  assign _zz_163 = _zz_130[32];
  assign _zz_164 = _zz_130[33];
  assign _zz_165 = _zz_130[34];
  assign _zz_166 = _zz_130[35];
  assign _zz_167 = _zz_130[36];
  assign _zz_168 = _zz_130[37];
  assign _zz_169 = _zz_130[38];
  assign _zz_170 = _zz_130[39];
  assign _zz_171 = _zz_130[40];
  assign _zz_172 = _zz_130[41];
  assign _zz_173 = _zz_130[42];
  assign _zz_174 = _zz_130[43];
  assign _zz_175 = _zz_130[44];
  assign _zz_176 = _zz_130[45];
  assign _zz_177 = _zz_130[46];
  assign _zz_178 = _zz_130[47];
  assign _zz_179 = _zz_130[48];
  assign _zz_180 = _zz_130[49];
  assign _zz_181 = _zz_130[50];
  assign _zz_182 = _zz_130[51];
  assign _zz_183 = _zz_130[52];
  assign _zz_184 = _zz_130[53];
  assign _zz_185 = _zz_130[54];
  assign _zz_186 = _zz_130[55];
  assign _zz_187 = _zz_130[56];
  assign _zz_188 = _zz_130[57];
  assign _zz_189 = _zz_130[58];
  assign _zz_190 = _zz_130[59];
  assign _zz_191 = _zz_130[60];
  assign _zz_192 = _zz_130[61];
  assign _zz_193 = _zz_130[62];
  assign _zz_194 = _zz_130[63];
  assign _zz_195 = _zz_130[64];
  assign _zz_196 = _zz_130[65];
  assign _zz_197 = _zz_130[66];
  assign _zz_198 = _zz_130[67];
  assign _zz_199 = _zz_130[68];
  assign _zz_200 = _zz_130[69];
  assign _zz_201 = _zz_130[70];
  assign _zz_202 = _zz_130[71];
  assign _zz_203 = _zz_130[72];
  assign _zz_204 = _zz_130[73];
  assign _zz_205 = _zz_130[74];
  assign _zz_206 = _zz_130[75];
  assign _zz_207 = _zz_130[76];
  assign _zz_208 = _zz_130[77];
  assign _zz_209 = _zz_130[78];
  assign _zz_210 = _zz_130[79];
  assign _zz_211 = _zz_130[80];
  assign _zz_212 = _zz_130[81];
  assign _zz_213 = _zz_130[82];
  assign _zz_214 = _zz_130[83];
  assign _zz_215 = _zz_130[84];
  assign _zz_216 = _zz_130[85];
  assign _zz_217 = _zz_130[86];
  assign _zz_218 = _zz_130[87];
  assign _zz_219 = _zz_130[88];
  assign _zz_220 = _zz_130[89];
  assign _zz_221 = _zz_130[90];
  assign _zz_222 = _zz_130[91];
  assign _zz_223 = _zz_130[92];
  assign _zz_224 = _zz_130[93];
  assign _zz_225 = _zz_130[94];
  assign _zz_226 = _zz_130[95];
  assign _zz_227 = _zz_130[96];
  assign _zz_228 = _zz_130[97];
  assign _zz_229 = _zz_130[98];
  assign _zz_230 = _zz_130[99];
  assign _zz_231 = _zz_130[100];
  assign _zz_232 = _zz_130[101];
  assign _zz_233 = _zz_130[102];
  assign _zz_234 = _zz_130[103];
  assign _zz_235 = _zz_130[104];
  assign _zz_236 = _zz_130[105];
  assign _zz_237 = _zz_130[106];
  assign _zz_238 = _zz_130[107];
  assign _zz_239 = _zz_130[108];
  assign _zz_240 = _zz_130[109];
  assign _zz_241 = _zz_130[110];
  assign _zz_242 = _zz_130[111];
  assign _zz_243 = _zz_130[112];
  assign _zz_244 = _zz_130[113];
  assign _zz_245 = _zz_130[114];
  assign _zz_246 = _zz_130[115];
  assign _zz_247 = _zz_130[116];
  assign _zz_248 = _zz_130[117];
  assign _zz_249 = _zz_130[118];
  assign _zz_250 = _zz_130[119];
  assign _zz_251 = _zz_130[120];
  assign _zz_252 = _zz_130[121];
  assign _zz_253 = _zz_130[122];
  assign _zz_254 = _zz_130[123];
  assign _zz_255 = _zz_130[124];
  assign _zz_256 = _zz_130[125];
  assign _zz_257 = _zz_130[126];
  assign _zz_258 = _zz_130[127];
  assign when_DCache_l217 = (is_hit && mru_full);
  assign when_DCache_l224 = (is_hit && cache_hit_0);
  assign when_DCache_l227 = (next_level_rdone && (2'b00 == evict_id_miss));
  assign when_DCache_l232 = (next_level_rdone && (2'b00 == evict_id_miss));
  assign when_DCache_l237 = ((flush || is_miss) || is_write);
  assign when_DCache_l240 = ((flush_done || next_level_rdone) || next_level_wdone);
  assign _zz_cache_hit_1 = _zz__zz_cache_hit_1;
  assign _zz_cache_mru_1 = _zz__zz_cache_mru_1;
  assign _zz_259 = ({127'd0,1'b1} <<< cpu_set);
  assign _zz_260 = _zz_259[0];
  assign _zz_261 = _zz_259[1];
  assign _zz_262 = _zz_259[2];
  assign _zz_263 = _zz_259[3];
  assign _zz_264 = _zz_259[4];
  assign _zz_265 = _zz_259[5];
  assign _zz_266 = _zz_259[6];
  assign _zz_267 = _zz_259[7];
  assign _zz_268 = _zz_259[8];
  assign _zz_269 = _zz_259[9];
  assign _zz_270 = _zz_259[10];
  assign _zz_271 = _zz_259[11];
  assign _zz_272 = _zz_259[12];
  assign _zz_273 = _zz_259[13];
  assign _zz_274 = _zz_259[14];
  assign _zz_275 = _zz_259[15];
  assign _zz_276 = _zz_259[16];
  assign _zz_277 = _zz_259[17];
  assign _zz_278 = _zz_259[18];
  assign _zz_279 = _zz_259[19];
  assign _zz_280 = _zz_259[20];
  assign _zz_281 = _zz_259[21];
  assign _zz_282 = _zz_259[22];
  assign _zz_283 = _zz_259[23];
  assign _zz_284 = _zz_259[24];
  assign _zz_285 = _zz_259[25];
  assign _zz_286 = _zz_259[26];
  assign _zz_287 = _zz_259[27];
  assign _zz_288 = _zz_259[28];
  assign _zz_289 = _zz_259[29];
  assign _zz_290 = _zz_259[30];
  assign _zz_291 = _zz_259[31];
  assign _zz_292 = _zz_259[32];
  assign _zz_293 = _zz_259[33];
  assign _zz_294 = _zz_259[34];
  assign _zz_295 = _zz_259[35];
  assign _zz_296 = _zz_259[36];
  assign _zz_297 = _zz_259[37];
  assign _zz_298 = _zz_259[38];
  assign _zz_299 = _zz_259[39];
  assign _zz_300 = _zz_259[40];
  assign _zz_301 = _zz_259[41];
  assign _zz_302 = _zz_259[42];
  assign _zz_303 = _zz_259[43];
  assign _zz_304 = _zz_259[44];
  assign _zz_305 = _zz_259[45];
  assign _zz_306 = _zz_259[46];
  assign _zz_307 = _zz_259[47];
  assign _zz_308 = _zz_259[48];
  assign _zz_309 = _zz_259[49];
  assign _zz_310 = _zz_259[50];
  assign _zz_311 = _zz_259[51];
  assign _zz_312 = _zz_259[52];
  assign _zz_313 = _zz_259[53];
  assign _zz_314 = _zz_259[54];
  assign _zz_315 = _zz_259[55];
  assign _zz_316 = _zz_259[56];
  assign _zz_317 = _zz_259[57];
  assign _zz_318 = _zz_259[58];
  assign _zz_319 = _zz_259[59];
  assign _zz_320 = _zz_259[60];
  assign _zz_321 = _zz_259[61];
  assign _zz_322 = _zz_259[62];
  assign _zz_323 = _zz_259[63];
  assign _zz_324 = _zz_259[64];
  assign _zz_325 = _zz_259[65];
  assign _zz_326 = _zz_259[66];
  assign _zz_327 = _zz_259[67];
  assign _zz_328 = _zz_259[68];
  assign _zz_329 = _zz_259[69];
  assign _zz_330 = _zz_259[70];
  assign _zz_331 = _zz_259[71];
  assign _zz_332 = _zz_259[72];
  assign _zz_333 = _zz_259[73];
  assign _zz_334 = _zz_259[74];
  assign _zz_335 = _zz_259[75];
  assign _zz_336 = _zz_259[76];
  assign _zz_337 = _zz_259[77];
  assign _zz_338 = _zz_259[78];
  assign _zz_339 = _zz_259[79];
  assign _zz_340 = _zz_259[80];
  assign _zz_341 = _zz_259[81];
  assign _zz_342 = _zz_259[82];
  assign _zz_343 = _zz_259[83];
  assign _zz_344 = _zz_259[84];
  assign _zz_345 = _zz_259[85];
  assign _zz_346 = _zz_259[86];
  assign _zz_347 = _zz_259[87];
  assign _zz_348 = _zz_259[88];
  assign _zz_349 = _zz_259[89];
  assign _zz_350 = _zz_259[90];
  assign _zz_351 = _zz_259[91];
  assign _zz_352 = _zz_259[92];
  assign _zz_353 = _zz_259[93];
  assign _zz_354 = _zz_259[94];
  assign _zz_355 = _zz_259[95];
  assign _zz_356 = _zz_259[96];
  assign _zz_357 = _zz_259[97];
  assign _zz_358 = _zz_259[98];
  assign _zz_359 = _zz_259[99];
  assign _zz_360 = _zz_259[100];
  assign _zz_361 = _zz_259[101];
  assign _zz_362 = _zz_259[102];
  assign _zz_363 = _zz_259[103];
  assign _zz_364 = _zz_259[104];
  assign _zz_365 = _zz_259[105];
  assign _zz_366 = _zz_259[106];
  assign _zz_367 = _zz_259[107];
  assign _zz_368 = _zz_259[108];
  assign _zz_369 = _zz_259[109];
  assign _zz_370 = _zz_259[110];
  assign _zz_371 = _zz_259[111];
  assign _zz_372 = _zz_259[112];
  assign _zz_373 = _zz_259[113];
  assign _zz_374 = _zz_259[114];
  assign _zz_375 = _zz_259[115];
  assign _zz_376 = _zz_259[116];
  assign _zz_377 = _zz_259[117];
  assign _zz_378 = _zz_259[118];
  assign _zz_379 = _zz_259[119];
  assign _zz_380 = _zz_259[120];
  assign _zz_381 = _zz_259[121];
  assign _zz_382 = _zz_259[122];
  assign _zz_383 = _zz_259[123];
  assign _zz_384 = _zz_259[124];
  assign _zz_385 = _zz_259[125];
  assign _zz_386 = _zz_259[126];
  assign _zz_387 = _zz_259[127];
  assign cache_tag_1 = _zz_cache_tag_1;
  assign cache_hit_1 = ((cache_tag_1 == cpu_tag) && _zz_cache_hit_1);
  assign cache_mru_1 = _zz_cache_mru_1;
  assign cache_invld_1 = (! _zz_cache_hit_1);
  assign cache_lru_1 = (! _zz_cache_mru_1);
  assign cache_victim_1 = (cache_invld_1 && cache_lru_1);
  assign sram_banks_data_1 = sram_1_ports_rsp_payload_data;
  assign sram_banks_valid_1 = sram_1_ports_rsp_valid;
  assign when_DCache_l181_1 = (is_hit && (2'b01 == hit_id));
  always @(*) begin
    if(when_DCache_l181_1) begin
      sram_1_ports_cmd_payload_addr = cpu_bank_addr;
    end else begin
      if(when_DCache_l188_1) begin
        sram_1_ports_cmd_payload_addr = cpu_bank_addr;
      end else begin
        if(when_DCache_l195_1) begin
          sram_1_ports_cmd_payload_addr = next_level_bank_addr;
        end else begin
          sram_1_ports_cmd_payload_addr = 7'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l181_1) begin
      sram_1_ports_cmd_valid = 1'b1;
    end else begin
      if(when_DCache_l188_1) begin
        sram_1_ports_cmd_valid = 1'b1;
      end else begin
        if(when_DCache_l195_1) begin
          sram_1_ports_cmd_valid = 1'b1;
        end else begin
          sram_1_ports_cmd_valid = 1'b0;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l181_1) begin
      sram_1_ports_cmd_payload_wen = ({7'h0,cpu_cmd_payload_wen} <<< cpu_bank_index);
    end else begin
      if(when_DCache_l188_1) begin
        sram_1_ports_cmd_payload_wen = 8'h0;
      end else begin
        if(when_DCache_l195_1) begin
          sram_1_ports_cmd_payload_wen = (_zz_sram_1_ports_cmd_payload_wen <<< _zz_sram_1_ports_cmd_payload_wen_1);
        end else begin
          sram_1_ports_cmd_payload_wen = 8'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l181_1) begin
      sram_1_ports_cmd_payload_wdata = ({448'h0,cpu_cmd_payload_wdata} <<< _zz_sram_1_ports_cmd_payload_wdata);
    end else begin
      if(when_DCache_l188_1) begin
        sram_1_ports_cmd_payload_wdata = 512'h0;
      end else begin
        if(when_DCache_l195_1) begin
          sram_1_ports_cmd_payload_wdata = ({448'h0,next_level_rsp_payload_data} <<< _zz_sram_1_ports_cmd_payload_wdata_1);
        end else begin
          sram_1_ports_cmd_payload_wdata = 512'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l181_1) begin
      sram_1_ports_cmd_payload_wstrb = ({56'h0,cpu_cmd_payload_wstrb} <<< _zz_sram_1_ports_cmd_payload_wstrb);
    end else begin
      if(when_DCache_l188_1) begin
        sram_1_ports_cmd_payload_wstrb = 64'h0;
      end else begin
        if(when_DCache_l195_1) begin
          sram_1_ports_cmd_payload_wstrb = ({56'h0,8'hff} <<< _zz_sram_1_ports_cmd_payload_wstrb_2);
        end else begin
          sram_1_ports_cmd_payload_wstrb = 64'h0;
        end
      end
    end
  end

  assign _zz_1034 = zz__zz_sram_1_ports_cmd_payload_wen(1'b0);
  always @(*) _zz_sram_1_ports_cmd_payload_wen = _zz_1034;
  assign when_DCache_l188_1 = ((next_level_rdone && (! is_write)) && (2'b01 == evict_id_miss));
  assign when_DCache_l195_1 = (next_level_rvalid && (2'b01 == evict_id_miss));
  assign _zz_388 = ({127'd0,1'b1} <<< flush_cnt_value);
  assign _zz_389 = _zz_388[0];
  assign _zz_390 = _zz_388[1];
  assign _zz_391 = _zz_388[2];
  assign _zz_392 = _zz_388[3];
  assign _zz_393 = _zz_388[4];
  assign _zz_394 = _zz_388[5];
  assign _zz_395 = _zz_388[6];
  assign _zz_396 = _zz_388[7];
  assign _zz_397 = _zz_388[8];
  assign _zz_398 = _zz_388[9];
  assign _zz_399 = _zz_388[10];
  assign _zz_400 = _zz_388[11];
  assign _zz_401 = _zz_388[12];
  assign _zz_402 = _zz_388[13];
  assign _zz_403 = _zz_388[14];
  assign _zz_404 = _zz_388[15];
  assign _zz_405 = _zz_388[16];
  assign _zz_406 = _zz_388[17];
  assign _zz_407 = _zz_388[18];
  assign _zz_408 = _zz_388[19];
  assign _zz_409 = _zz_388[20];
  assign _zz_410 = _zz_388[21];
  assign _zz_411 = _zz_388[22];
  assign _zz_412 = _zz_388[23];
  assign _zz_413 = _zz_388[24];
  assign _zz_414 = _zz_388[25];
  assign _zz_415 = _zz_388[26];
  assign _zz_416 = _zz_388[27];
  assign _zz_417 = _zz_388[28];
  assign _zz_418 = _zz_388[29];
  assign _zz_419 = _zz_388[30];
  assign _zz_420 = _zz_388[31];
  assign _zz_421 = _zz_388[32];
  assign _zz_422 = _zz_388[33];
  assign _zz_423 = _zz_388[34];
  assign _zz_424 = _zz_388[35];
  assign _zz_425 = _zz_388[36];
  assign _zz_426 = _zz_388[37];
  assign _zz_427 = _zz_388[38];
  assign _zz_428 = _zz_388[39];
  assign _zz_429 = _zz_388[40];
  assign _zz_430 = _zz_388[41];
  assign _zz_431 = _zz_388[42];
  assign _zz_432 = _zz_388[43];
  assign _zz_433 = _zz_388[44];
  assign _zz_434 = _zz_388[45];
  assign _zz_435 = _zz_388[46];
  assign _zz_436 = _zz_388[47];
  assign _zz_437 = _zz_388[48];
  assign _zz_438 = _zz_388[49];
  assign _zz_439 = _zz_388[50];
  assign _zz_440 = _zz_388[51];
  assign _zz_441 = _zz_388[52];
  assign _zz_442 = _zz_388[53];
  assign _zz_443 = _zz_388[54];
  assign _zz_444 = _zz_388[55];
  assign _zz_445 = _zz_388[56];
  assign _zz_446 = _zz_388[57];
  assign _zz_447 = _zz_388[58];
  assign _zz_448 = _zz_388[59];
  assign _zz_449 = _zz_388[60];
  assign _zz_450 = _zz_388[61];
  assign _zz_451 = _zz_388[62];
  assign _zz_452 = _zz_388[63];
  assign _zz_453 = _zz_388[64];
  assign _zz_454 = _zz_388[65];
  assign _zz_455 = _zz_388[66];
  assign _zz_456 = _zz_388[67];
  assign _zz_457 = _zz_388[68];
  assign _zz_458 = _zz_388[69];
  assign _zz_459 = _zz_388[70];
  assign _zz_460 = _zz_388[71];
  assign _zz_461 = _zz_388[72];
  assign _zz_462 = _zz_388[73];
  assign _zz_463 = _zz_388[74];
  assign _zz_464 = _zz_388[75];
  assign _zz_465 = _zz_388[76];
  assign _zz_466 = _zz_388[77];
  assign _zz_467 = _zz_388[78];
  assign _zz_468 = _zz_388[79];
  assign _zz_469 = _zz_388[80];
  assign _zz_470 = _zz_388[81];
  assign _zz_471 = _zz_388[82];
  assign _zz_472 = _zz_388[83];
  assign _zz_473 = _zz_388[84];
  assign _zz_474 = _zz_388[85];
  assign _zz_475 = _zz_388[86];
  assign _zz_476 = _zz_388[87];
  assign _zz_477 = _zz_388[88];
  assign _zz_478 = _zz_388[89];
  assign _zz_479 = _zz_388[90];
  assign _zz_480 = _zz_388[91];
  assign _zz_481 = _zz_388[92];
  assign _zz_482 = _zz_388[93];
  assign _zz_483 = _zz_388[94];
  assign _zz_484 = _zz_388[95];
  assign _zz_485 = _zz_388[96];
  assign _zz_486 = _zz_388[97];
  assign _zz_487 = _zz_388[98];
  assign _zz_488 = _zz_388[99];
  assign _zz_489 = _zz_388[100];
  assign _zz_490 = _zz_388[101];
  assign _zz_491 = _zz_388[102];
  assign _zz_492 = _zz_388[103];
  assign _zz_493 = _zz_388[104];
  assign _zz_494 = _zz_388[105];
  assign _zz_495 = _zz_388[106];
  assign _zz_496 = _zz_388[107];
  assign _zz_497 = _zz_388[108];
  assign _zz_498 = _zz_388[109];
  assign _zz_499 = _zz_388[110];
  assign _zz_500 = _zz_388[111];
  assign _zz_501 = _zz_388[112];
  assign _zz_502 = _zz_388[113];
  assign _zz_503 = _zz_388[114];
  assign _zz_504 = _zz_388[115];
  assign _zz_505 = _zz_388[116];
  assign _zz_506 = _zz_388[117];
  assign _zz_507 = _zz_388[118];
  assign _zz_508 = _zz_388[119];
  assign _zz_509 = _zz_388[120];
  assign _zz_510 = _zz_388[121];
  assign _zz_511 = _zz_388[122];
  assign _zz_512 = _zz_388[123];
  assign _zz_513 = _zz_388[124];
  assign _zz_514 = _zz_388[125];
  assign _zz_515 = _zz_388[126];
  assign _zz_516 = _zz_388[127];
  assign when_DCache_l217_1 = (is_hit && mru_full);
  assign when_DCache_l224_1 = (is_hit && cache_hit_1);
  assign when_DCache_l227_1 = (next_level_rdone && (2'b01 == evict_id_miss));
  assign when_DCache_l232_1 = (next_level_rdone && (2'b01 == evict_id_miss));
  assign when_DCache_l237_1 = ((flush || is_miss) || is_write);
  assign when_DCache_l240_1 = ((flush_done || next_level_rdone) || next_level_wdone);
  assign _zz_cache_hit_2 = _zz__zz_cache_hit_2;
  assign _zz_cache_mru_2 = _zz__zz_cache_mru_2;
  assign _zz_517 = ({127'd0,1'b1} <<< cpu_set);
  assign _zz_518 = _zz_517[0];
  assign _zz_519 = _zz_517[1];
  assign _zz_520 = _zz_517[2];
  assign _zz_521 = _zz_517[3];
  assign _zz_522 = _zz_517[4];
  assign _zz_523 = _zz_517[5];
  assign _zz_524 = _zz_517[6];
  assign _zz_525 = _zz_517[7];
  assign _zz_526 = _zz_517[8];
  assign _zz_527 = _zz_517[9];
  assign _zz_528 = _zz_517[10];
  assign _zz_529 = _zz_517[11];
  assign _zz_530 = _zz_517[12];
  assign _zz_531 = _zz_517[13];
  assign _zz_532 = _zz_517[14];
  assign _zz_533 = _zz_517[15];
  assign _zz_534 = _zz_517[16];
  assign _zz_535 = _zz_517[17];
  assign _zz_536 = _zz_517[18];
  assign _zz_537 = _zz_517[19];
  assign _zz_538 = _zz_517[20];
  assign _zz_539 = _zz_517[21];
  assign _zz_540 = _zz_517[22];
  assign _zz_541 = _zz_517[23];
  assign _zz_542 = _zz_517[24];
  assign _zz_543 = _zz_517[25];
  assign _zz_544 = _zz_517[26];
  assign _zz_545 = _zz_517[27];
  assign _zz_546 = _zz_517[28];
  assign _zz_547 = _zz_517[29];
  assign _zz_548 = _zz_517[30];
  assign _zz_549 = _zz_517[31];
  assign _zz_550 = _zz_517[32];
  assign _zz_551 = _zz_517[33];
  assign _zz_552 = _zz_517[34];
  assign _zz_553 = _zz_517[35];
  assign _zz_554 = _zz_517[36];
  assign _zz_555 = _zz_517[37];
  assign _zz_556 = _zz_517[38];
  assign _zz_557 = _zz_517[39];
  assign _zz_558 = _zz_517[40];
  assign _zz_559 = _zz_517[41];
  assign _zz_560 = _zz_517[42];
  assign _zz_561 = _zz_517[43];
  assign _zz_562 = _zz_517[44];
  assign _zz_563 = _zz_517[45];
  assign _zz_564 = _zz_517[46];
  assign _zz_565 = _zz_517[47];
  assign _zz_566 = _zz_517[48];
  assign _zz_567 = _zz_517[49];
  assign _zz_568 = _zz_517[50];
  assign _zz_569 = _zz_517[51];
  assign _zz_570 = _zz_517[52];
  assign _zz_571 = _zz_517[53];
  assign _zz_572 = _zz_517[54];
  assign _zz_573 = _zz_517[55];
  assign _zz_574 = _zz_517[56];
  assign _zz_575 = _zz_517[57];
  assign _zz_576 = _zz_517[58];
  assign _zz_577 = _zz_517[59];
  assign _zz_578 = _zz_517[60];
  assign _zz_579 = _zz_517[61];
  assign _zz_580 = _zz_517[62];
  assign _zz_581 = _zz_517[63];
  assign _zz_582 = _zz_517[64];
  assign _zz_583 = _zz_517[65];
  assign _zz_584 = _zz_517[66];
  assign _zz_585 = _zz_517[67];
  assign _zz_586 = _zz_517[68];
  assign _zz_587 = _zz_517[69];
  assign _zz_588 = _zz_517[70];
  assign _zz_589 = _zz_517[71];
  assign _zz_590 = _zz_517[72];
  assign _zz_591 = _zz_517[73];
  assign _zz_592 = _zz_517[74];
  assign _zz_593 = _zz_517[75];
  assign _zz_594 = _zz_517[76];
  assign _zz_595 = _zz_517[77];
  assign _zz_596 = _zz_517[78];
  assign _zz_597 = _zz_517[79];
  assign _zz_598 = _zz_517[80];
  assign _zz_599 = _zz_517[81];
  assign _zz_600 = _zz_517[82];
  assign _zz_601 = _zz_517[83];
  assign _zz_602 = _zz_517[84];
  assign _zz_603 = _zz_517[85];
  assign _zz_604 = _zz_517[86];
  assign _zz_605 = _zz_517[87];
  assign _zz_606 = _zz_517[88];
  assign _zz_607 = _zz_517[89];
  assign _zz_608 = _zz_517[90];
  assign _zz_609 = _zz_517[91];
  assign _zz_610 = _zz_517[92];
  assign _zz_611 = _zz_517[93];
  assign _zz_612 = _zz_517[94];
  assign _zz_613 = _zz_517[95];
  assign _zz_614 = _zz_517[96];
  assign _zz_615 = _zz_517[97];
  assign _zz_616 = _zz_517[98];
  assign _zz_617 = _zz_517[99];
  assign _zz_618 = _zz_517[100];
  assign _zz_619 = _zz_517[101];
  assign _zz_620 = _zz_517[102];
  assign _zz_621 = _zz_517[103];
  assign _zz_622 = _zz_517[104];
  assign _zz_623 = _zz_517[105];
  assign _zz_624 = _zz_517[106];
  assign _zz_625 = _zz_517[107];
  assign _zz_626 = _zz_517[108];
  assign _zz_627 = _zz_517[109];
  assign _zz_628 = _zz_517[110];
  assign _zz_629 = _zz_517[111];
  assign _zz_630 = _zz_517[112];
  assign _zz_631 = _zz_517[113];
  assign _zz_632 = _zz_517[114];
  assign _zz_633 = _zz_517[115];
  assign _zz_634 = _zz_517[116];
  assign _zz_635 = _zz_517[117];
  assign _zz_636 = _zz_517[118];
  assign _zz_637 = _zz_517[119];
  assign _zz_638 = _zz_517[120];
  assign _zz_639 = _zz_517[121];
  assign _zz_640 = _zz_517[122];
  assign _zz_641 = _zz_517[123];
  assign _zz_642 = _zz_517[124];
  assign _zz_643 = _zz_517[125];
  assign _zz_644 = _zz_517[126];
  assign _zz_645 = _zz_517[127];
  assign cache_tag_2 = _zz_cache_tag_2;
  assign cache_hit_2 = ((cache_tag_2 == cpu_tag) && _zz_cache_hit_2);
  assign cache_mru_2 = _zz_cache_mru_2;
  assign cache_invld_2 = (! _zz_cache_hit_2);
  assign cache_lru_2 = (! _zz_cache_mru_2);
  assign cache_victim_2 = (cache_invld_2 && cache_lru_2);
  assign sram_banks_data_2 = sram_2_ports_rsp_payload_data;
  assign sram_banks_valid_2 = sram_2_ports_rsp_valid;
  assign when_DCache_l181_2 = (is_hit && (2'b10 == hit_id));
  always @(*) begin
    if(when_DCache_l181_2) begin
      sram_2_ports_cmd_payload_addr = cpu_bank_addr;
    end else begin
      if(when_DCache_l188_2) begin
        sram_2_ports_cmd_payload_addr = cpu_bank_addr;
      end else begin
        if(when_DCache_l195_2) begin
          sram_2_ports_cmd_payload_addr = next_level_bank_addr;
        end else begin
          sram_2_ports_cmd_payload_addr = 7'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l181_2) begin
      sram_2_ports_cmd_valid = 1'b1;
    end else begin
      if(when_DCache_l188_2) begin
        sram_2_ports_cmd_valid = 1'b1;
      end else begin
        if(when_DCache_l195_2) begin
          sram_2_ports_cmd_valid = 1'b1;
        end else begin
          sram_2_ports_cmd_valid = 1'b0;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l181_2) begin
      sram_2_ports_cmd_payload_wen = ({7'h0,cpu_cmd_payload_wen} <<< cpu_bank_index);
    end else begin
      if(when_DCache_l188_2) begin
        sram_2_ports_cmd_payload_wen = 8'h0;
      end else begin
        if(when_DCache_l195_2) begin
          sram_2_ports_cmd_payload_wen = (_zz_sram_2_ports_cmd_payload_wen <<< _zz_sram_2_ports_cmd_payload_wen_1);
        end else begin
          sram_2_ports_cmd_payload_wen = 8'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l181_2) begin
      sram_2_ports_cmd_payload_wdata = ({448'h0,cpu_cmd_payload_wdata} <<< _zz_sram_2_ports_cmd_payload_wdata);
    end else begin
      if(when_DCache_l188_2) begin
        sram_2_ports_cmd_payload_wdata = 512'h0;
      end else begin
        if(when_DCache_l195_2) begin
          sram_2_ports_cmd_payload_wdata = ({448'h0,next_level_rsp_payload_data} <<< _zz_sram_2_ports_cmd_payload_wdata_1);
        end else begin
          sram_2_ports_cmd_payload_wdata = 512'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l181_2) begin
      sram_2_ports_cmd_payload_wstrb = ({56'h0,cpu_cmd_payload_wstrb} <<< _zz_sram_2_ports_cmd_payload_wstrb);
    end else begin
      if(when_DCache_l188_2) begin
        sram_2_ports_cmd_payload_wstrb = 64'h0;
      end else begin
        if(when_DCache_l195_2) begin
          sram_2_ports_cmd_payload_wstrb = ({56'h0,8'hff} <<< _zz_sram_2_ports_cmd_payload_wstrb_2);
        end else begin
          sram_2_ports_cmd_payload_wstrb = 64'h0;
        end
      end
    end
  end

  assign _zz_1035 = zz__zz_sram_2_ports_cmd_payload_wen(1'b0);
  always @(*) _zz_sram_2_ports_cmd_payload_wen = _zz_1035;
  assign when_DCache_l188_2 = ((next_level_rdone && (! is_write)) && (2'b10 == evict_id_miss));
  assign when_DCache_l195_2 = (next_level_rvalid && (2'b10 == evict_id_miss));
  assign _zz_646 = ({127'd0,1'b1} <<< flush_cnt_value);
  assign _zz_647 = _zz_646[0];
  assign _zz_648 = _zz_646[1];
  assign _zz_649 = _zz_646[2];
  assign _zz_650 = _zz_646[3];
  assign _zz_651 = _zz_646[4];
  assign _zz_652 = _zz_646[5];
  assign _zz_653 = _zz_646[6];
  assign _zz_654 = _zz_646[7];
  assign _zz_655 = _zz_646[8];
  assign _zz_656 = _zz_646[9];
  assign _zz_657 = _zz_646[10];
  assign _zz_658 = _zz_646[11];
  assign _zz_659 = _zz_646[12];
  assign _zz_660 = _zz_646[13];
  assign _zz_661 = _zz_646[14];
  assign _zz_662 = _zz_646[15];
  assign _zz_663 = _zz_646[16];
  assign _zz_664 = _zz_646[17];
  assign _zz_665 = _zz_646[18];
  assign _zz_666 = _zz_646[19];
  assign _zz_667 = _zz_646[20];
  assign _zz_668 = _zz_646[21];
  assign _zz_669 = _zz_646[22];
  assign _zz_670 = _zz_646[23];
  assign _zz_671 = _zz_646[24];
  assign _zz_672 = _zz_646[25];
  assign _zz_673 = _zz_646[26];
  assign _zz_674 = _zz_646[27];
  assign _zz_675 = _zz_646[28];
  assign _zz_676 = _zz_646[29];
  assign _zz_677 = _zz_646[30];
  assign _zz_678 = _zz_646[31];
  assign _zz_679 = _zz_646[32];
  assign _zz_680 = _zz_646[33];
  assign _zz_681 = _zz_646[34];
  assign _zz_682 = _zz_646[35];
  assign _zz_683 = _zz_646[36];
  assign _zz_684 = _zz_646[37];
  assign _zz_685 = _zz_646[38];
  assign _zz_686 = _zz_646[39];
  assign _zz_687 = _zz_646[40];
  assign _zz_688 = _zz_646[41];
  assign _zz_689 = _zz_646[42];
  assign _zz_690 = _zz_646[43];
  assign _zz_691 = _zz_646[44];
  assign _zz_692 = _zz_646[45];
  assign _zz_693 = _zz_646[46];
  assign _zz_694 = _zz_646[47];
  assign _zz_695 = _zz_646[48];
  assign _zz_696 = _zz_646[49];
  assign _zz_697 = _zz_646[50];
  assign _zz_698 = _zz_646[51];
  assign _zz_699 = _zz_646[52];
  assign _zz_700 = _zz_646[53];
  assign _zz_701 = _zz_646[54];
  assign _zz_702 = _zz_646[55];
  assign _zz_703 = _zz_646[56];
  assign _zz_704 = _zz_646[57];
  assign _zz_705 = _zz_646[58];
  assign _zz_706 = _zz_646[59];
  assign _zz_707 = _zz_646[60];
  assign _zz_708 = _zz_646[61];
  assign _zz_709 = _zz_646[62];
  assign _zz_710 = _zz_646[63];
  assign _zz_711 = _zz_646[64];
  assign _zz_712 = _zz_646[65];
  assign _zz_713 = _zz_646[66];
  assign _zz_714 = _zz_646[67];
  assign _zz_715 = _zz_646[68];
  assign _zz_716 = _zz_646[69];
  assign _zz_717 = _zz_646[70];
  assign _zz_718 = _zz_646[71];
  assign _zz_719 = _zz_646[72];
  assign _zz_720 = _zz_646[73];
  assign _zz_721 = _zz_646[74];
  assign _zz_722 = _zz_646[75];
  assign _zz_723 = _zz_646[76];
  assign _zz_724 = _zz_646[77];
  assign _zz_725 = _zz_646[78];
  assign _zz_726 = _zz_646[79];
  assign _zz_727 = _zz_646[80];
  assign _zz_728 = _zz_646[81];
  assign _zz_729 = _zz_646[82];
  assign _zz_730 = _zz_646[83];
  assign _zz_731 = _zz_646[84];
  assign _zz_732 = _zz_646[85];
  assign _zz_733 = _zz_646[86];
  assign _zz_734 = _zz_646[87];
  assign _zz_735 = _zz_646[88];
  assign _zz_736 = _zz_646[89];
  assign _zz_737 = _zz_646[90];
  assign _zz_738 = _zz_646[91];
  assign _zz_739 = _zz_646[92];
  assign _zz_740 = _zz_646[93];
  assign _zz_741 = _zz_646[94];
  assign _zz_742 = _zz_646[95];
  assign _zz_743 = _zz_646[96];
  assign _zz_744 = _zz_646[97];
  assign _zz_745 = _zz_646[98];
  assign _zz_746 = _zz_646[99];
  assign _zz_747 = _zz_646[100];
  assign _zz_748 = _zz_646[101];
  assign _zz_749 = _zz_646[102];
  assign _zz_750 = _zz_646[103];
  assign _zz_751 = _zz_646[104];
  assign _zz_752 = _zz_646[105];
  assign _zz_753 = _zz_646[106];
  assign _zz_754 = _zz_646[107];
  assign _zz_755 = _zz_646[108];
  assign _zz_756 = _zz_646[109];
  assign _zz_757 = _zz_646[110];
  assign _zz_758 = _zz_646[111];
  assign _zz_759 = _zz_646[112];
  assign _zz_760 = _zz_646[113];
  assign _zz_761 = _zz_646[114];
  assign _zz_762 = _zz_646[115];
  assign _zz_763 = _zz_646[116];
  assign _zz_764 = _zz_646[117];
  assign _zz_765 = _zz_646[118];
  assign _zz_766 = _zz_646[119];
  assign _zz_767 = _zz_646[120];
  assign _zz_768 = _zz_646[121];
  assign _zz_769 = _zz_646[122];
  assign _zz_770 = _zz_646[123];
  assign _zz_771 = _zz_646[124];
  assign _zz_772 = _zz_646[125];
  assign _zz_773 = _zz_646[126];
  assign _zz_774 = _zz_646[127];
  assign when_DCache_l217_2 = (is_hit && mru_full);
  assign when_DCache_l224_2 = (is_hit && cache_hit_2);
  assign when_DCache_l227_2 = (next_level_rdone && (2'b10 == evict_id_miss));
  assign when_DCache_l232_2 = (next_level_rdone && (2'b10 == evict_id_miss));
  assign when_DCache_l237_2 = ((flush || is_miss) || is_write);
  assign when_DCache_l240_2 = ((flush_done || next_level_rdone) || next_level_wdone);
  assign _zz_cache_hit_3 = _zz__zz_cache_hit_3;
  assign _zz_cache_mru_3 = _zz__zz_cache_mru_3;
  assign _zz_775 = ({127'd0,1'b1} <<< cpu_set);
  assign _zz_776 = _zz_775[0];
  assign _zz_777 = _zz_775[1];
  assign _zz_778 = _zz_775[2];
  assign _zz_779 = _zz_775[3];
  assign _zz_780 = _zz_775[4];
  assign _zz_781 = _zz_775[5];
  assign _zz_782 = _zz_775[6];
  assign _zz_783 = _zz_775[7];
  assign _zz_784 = _zz_775[8];
  assign _zz_785 = _zz_775[9];
  assign _zz_786 = _zz_775[10];
  assign _zz_787 = _zz_775[11];
  assign _zz_788 = _zz_775[12];
  assign _zz_789 = _zz_775[13];
  assign _zz_790 = _zz_775[14];
  assign _zz_791 = _zz_775[15];
  assign _zz_792 = _zz_775[16];
  assign _zz_793 = _zz_775[17];
  assign _zz_794 = _zz_775[18];
  assign _zz_795 = _zz_775[19];
  assign _zz_796 = _zz_775[20];
  assign _zz_797 = _zz_775[21];
  assign _zz_798 = _zz_775[22];
  assign _zz_799 = _zz_775[23];
  assign _zz_800 = _zz_775[24];
  assign _zz_801 = _zz_775[25];
  assign _zz_802 = _zz_775[26];
  assign _zz_803 = _zz_775[27];
  assign _zz_804 = _zz_775[28];
  assign _zz_805 = _zz_775[29];
  assign _zz_806 = _zz_775[30];
  assign _zz_807 = _zz_775[31];
  assign _zz_808 = _zz_775[32];
  assign _zz_809 = _zz_775[33];
  assign _zz_810 = _zz_775[34];
  assign _zz_811 = _zz_775[35];
  assign _zz_812 = _zz_775[36];
  assign _zz_813 = _zz_775[37];
  assign _zz_814 = _zz_775[38];
  assign _zz_815 = _zz_775[39];
  assign _zz_816 = _zz_775[40];
  assign _zz_817 = _zz_775[41];
  assign _zz_818 = _zz_775[42];
  assign _zz_819 = _zz_775[43];
  assign _zz_820 = _zz_775[44];
  assign _zz_821 = _zz_775[45];
  assign _zz_822 = _zz_775[46];
  assign _zz_823 = _zz_775[47];
  assign _zz_824 = _zz_775[48];
  assign _zz_825 = _zz_775[49];
  assign _zz_826 = _zz_775[50];
  assign _zz_827 = _zz_775[51];
  assign _zz_828 = _zz_775[52];
  assign _zz_829 = _zz_775[53];
  assign _zz_830 = _zz_775[54];
  assign _zz_831 = _zz_775[55];
  assign _zz_832 = _zz_775[56];
  assign _zz_833 = _zz_775[57];
  assign _zz_834 = _zz_775[58];
  assign _zz_835 = _zz_775[59];
  assign _zz_836 = _zz_775[60];
  assign _zz_837 = _zz_775[61];
  assign _zz_838 = _zz_775[62];
  assign _zz_839 = _zz_775[63];
  assign _zz_840 = _zz_775[64];
  assign _zz_841 = _zz_775[65];
  assign _zz_842 = _zz_775[66];
  assign _zz_843 = _zz_775[67];
  assign _zz_844 = _zz_775[68];
  assign _zz_845 = _zz_775[69];
  assign _zz_846 = _zz_775[70];
  assign _zz_847 = _zz_775[71];
  assign _zz_848 = _zz_775[72];
  assign _zz_849 = _zz_775[73];
  assign _zz_850 = _zz_775[74];
  assign _zz_851 = _zz_775[75];
  assign _zz_852 = _zz_775[76];
  assign _zz_853 = _zz_775[77];
  assign _zz_854 = _zz_775[78];
  assign _zz_855 = _zz_775[79];
  assign _zz_856 = _zz_775[80];
  assign _zz_857 = _zz_775[81];
  assign _zz_858 = _zz_775[82];
  assign _zz_859 = _zz_775[83];
  assign _zz_860 = _zz_775[84];
  assign _zz_861 = _zz_775[85];
  assign _zz_862 = _zz_775[86];
  assign _zz_863 = _zz_775[87];
  assign _zz_864 = _zz_775[88];
  assign _zz_865 = _zz_775[89];
  assign _zz_866 = _zz_775[90];
  assign _zz_867 = _zz_775[91];
  assign _zz_868 = _zz_775[92];
  assign _zz_869 = _zz_775[93];
  assign _zz_870 = _zz_775[94];
  assign _zz_871 = _zz_775[95];
  assign _zz_872 = _zz_775[96];
  assign _zz_873 = _zz_775[97];
  assign _zz_874 = _zz_775[98];
  assign _zz_875 = _zz_775[99];
  assign _zz_876 = _zz_775[100];
  assign _zz_877 = _zz_775[101];
  assign _zz_878 = _zz_775[102];
  assign _zz_879 = _zz_775[103];
  assign _zz_880 = _zz_775[104];
  assign _zz_881 = _zz_775[105];
  assign _zz_882 = _zz_775[106];
  assign _zz_883 = _zz_775[107];
  assign _zz_884 = _zz_775[108];
  assign _zz_885 = _zz_775[109];
  assign _zz_886 = _zz_775[110];
  assign _zz_887 = _zz_775[111];
  assign _zz_888 = _zz_775[112];
  assign _zz_889 = _zz_775[113];
  assign _zz_890 = _zz_775[114];
  assign _zz_891 = _zz_775[115];
  assign _zz_892 = _zz_775[116];
  assign _zz_893 = _zz_775[117];
  assign _zz_894 = _zz_775[118];
  assign _zz_895 = _zz_775[119];
  assign _zz_896 = _zz_775[120];
  assign _zz_897 = _zz_775[121];
  assign _zz_898 = _zz_775[122];
  assign _zz_899 = _zz_775[123];
  assign _zz_900 = _zz_775[124];
  assign _zz_901 = _zz_775[125];
  assign _zz_902 = _zz_775[126];
  assign _zz_903 = _zz_775[127];
  assign cache_tag_3 = _zz_cache_tag_3;
  assign cache_hit_3 = ((cache_tag_3 == cpu_tag) && _zz_cache_hit_3);
  assign cache_mru_3 = _zz_cache_mru_3;
  assign cache_invld_3 = (! _zz_cache_hit_3);
  assign cache_lru_3 = (! _zz_cache_mru_3);
  assign cache_victim_3 = (cache_invld_3 && cache_lru_3);
  assign sram_banks_data_3 = sram_3_ports_rsp_payload_data;
  assign sram_banks_valid_3 = sram_3_ports_rsp_valid;
  assign when_DCache_l181_3 = (is_hit && (2'b11 == hit_id));
  always @(*) begin
    if(when_DCache_l181_3) begin
      sram_3_ports_cmd_payload_addr = cpu_bank_addr;
    end else begin
      if(when_DCache_l188_3) begin
        sram_3_ports_cmd_payload_addr = cpu_bank_addr;
      end else begin
        if(when_DCache_l195_3) begin
          sram_3_ports_cmd_payload_addr = next_level_bank_addr;
        end else begin
          sram_3_ports_cmd_payload_addr = 7'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l181_3) begin
      sram_3_ports_cmd_valid = 1'b1;
    end else begin
      if(when_DCache_l188_3) begin
        sram_3_ports_cmd_valid = 1'b1;
      end else begin
        if(when_DCache_l195_3) begin
          sram_3_ports_cmd_valid = 1'b1;
        end else begin
          sram_3_ports_cmd_valid = 1'b0;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l181_3) begin
      sram_3_ports_cmd_payload_wen = ({7'h0,cpu_cmd_payload_wen} <<< cpu_bank_index);
    end else begin
      if(when_DCache_l188_3) begin
        sram_3_ports_cmd_payload_wen = 8'h0;
      end else begin
        if(when_DCache_l195_3) begin
          sram_3_ports_cmd_payload_wen = (_zz_sram_3_ports_cmd_payload_wen <<< _zz_sram_3_ports_cmd_payload_wen_1);
        end else begin
          sram_3_ports_cmd_payload_wen = 8'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l181_3) begin
      sram_3_ports_cmd_payload_wdata = ({448'h0,cpu_cmd_payload_wdata} <<< _zz_sram_3_ports_cmd_payload_wdata);
    end else begin
      if(when_DCache_l188_3) begin
        sram_3_ports_cmd_payload_wdata = 512'h0;
      end else begin
        if(when_DCache_l195_3) begin
          sram_3_ports_cmd_payload_wdata = ({448'h0,next_level_rsp_payload_data} <<< _zz_sram_3_ports_cmd_payload_wdata_1);
        end else begin
          sram_3_ports_cmd_payload_wdata = 512'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_DCache_l181_3) begin
      sram_3_ports_cmd_payload_wstrb = ({56'h0,cpu_cmd_payload_wstrb} <<< _zz_sram_3_ports_cmd_payload_wstrb);
    end else begin
      if(when_DCache_l188_3) begin
        sram_3_ports_cmd_payload_wstrb = 64'h0;
      end else begin
        if(when_DCache_l195_3) begin
          sram_3_ports_cmd_payload_wstrb = ({56'h0,8'hff} <<< _zz_sram_3_ports_cmd_payload_wstrb_2);
        end else begin
          sram_3_ports_cmd_payload_wstrb = 64'h0;
        end
      end
    end
  end

  assign _zz_1036 = zz__zz_sram_3_ports_cmd_payload_wen(1'b0);
  always @(*) _zz_sram_3_ports_cmd_payload_wen = _zz_1036;
  assign when_DCache_l188_3 = ((next_level_rdone && (! is_write)) && (2'b11 == evict_id_miss));
  assign when_DCache_l195_3 = (next_level_rvalid && (2'b11 == evict_id_miss));
  assign _zz_904 = ({127'd0,1'b1} <<< flush_cnt_value);
  assign _zz_905 = _zz_904[0];
  assign _zz_906 = _zz_904[1];
  assign _zz_907 = _zz_904[2];
  assign _zz_908 = _zz_904[3];
  assign _zz_909 = _zz_904[4];
  assign _zz_910 = _zz_904[5];
  assign _zz_911 = _zz_904[6];
  assign _zz_912 = _zz_904[7];
  assign _zz_913 = _zz_904[8];
  assign _zz_914 = _zz_904[9];
  assign _zz_915 = _zz_904[10];
  assign _zz_916 = _zz_904[11];
  assign _zz_917 = _zz_904[12];
  assign _zz_918 = _zz_904[13];
  assign _zz_919 = _zz_904[14];
  assign _zz_920 = _zz_904[15];
  assign _zz_921 = _zz_904[16];
  assign _zz_922 = _zz_904[17];
  assign _zz_923 = _zz_904[18];
  assign _zz_924 = _zz_904[19];
  assign _zz_925 = _zz_904[20];
  assign _zz_926 = _zz_904[21];
  assign _zz_927 = _zz_904[22];
  assign _zz_928 = _zz_904[23];
  assign _zz_929 = _zz_904[24];
  assign _zz_930 = _zz_904[25];
  assign _zz_931 = _zz_904[26];
  assign _zz_932 = _zz_904[27];
  assign _zz_933 = _zz_904[28];
  assign _zz_934 = _zz_904[29];
  assign _zz_935 = _zz_904[30];
  assign _zz_936 = _zz_904[31];
  assign _zz_937 = _zz_904[32];
  assign _zz_938 = _zz_904[33];
  assign _zz_939 = _zz_904[34];
  assign _zz_940 = _zz_904[35];
  assign _zz_941 = _zz_904[36];
  assign _zz_942 = _zz_904[37];
  assign _zz_943 = _zz_904[38];
  assign _zz_944 = _zz_904[39];
  assign _zz_945 = _zz_904[40];
  assign _zz_946 = _zz_904[41];
  assign _zz_947 = _zz_904[42];
  assign _zz_948 = _zz_904[43];
  assign _zz_949 = _zz_904[44];
  assign _zz_950 = _zz_904[45];
  assign _zz_951 = _zz_904[46];
  assign _zz_952 = _zz_904[47];
  assign _zz_953 = _zz_904[48];
  assign _zz_954 = _zz_904[49];
  assign _zz_955 = _zz_904[50];
  assign _zz_956 = _zz_904[51];
  assign _zz_957 = _zz_904[52];
  assign _zz_958 = _zz_904[53];
  assign _zz_959 = _zz_904[54];
  assign _zz_960 = _zz_904[55];
  assign _zz_961 = _zz_904[56];
  assign _zz_962 = _zz_904[57];
  assign _zz_963 = _zz_904[58];
  assign _zz_964 = _zz_904[59];
  assign _zz_965 = _zz_904[60];
  assign _zz_966 = _zz_904[61];
  assign _zz_967 = _zz_904[62];
  assign _zz_968 = _zz_904[63];
  assign _zz_969 = _zz_904[64];
  assign _zz_970 = _zz_904[65];
  assign _zz_971 = _zz_904[66];
  assign _zz_972 = _zz_904[67];
  assign _zz_973 = _zz_904[68];
  assign _zz_974 = _zz_904[69];
  assign _zz_975 = _zz_904[70];
  assign _zz_976 = _zz_904[71];
  assign _zz_977 = _zz_904[72];
  assign _zz_978 = _zz_904[73];
  assign _zz_979 = _zz_904[74];
  assign _zz_980 = _zz_904[75];
  assign _zz_981 = _zz_904[76];
  assign _zz_982 = _zz_904[77];
  assign _zz_983 = _zz_904[78];
  assign _zz_984 = _zz_904[79];
  assign _zz_985 = _zz_904[80];
  assign _zz_986 = _zz_904[81];
  assign _zz_987 = _zz_904[82];
  assign _zz_988 = _zz_904[83];
  assign _zz_989 = _zz_904[84];
  assign _zz_990 = _zz_904[85];
  assign _zz_991 = _zz_904[86];
  assign _zz_992 = _zz_904[87];
  assign _zz_993 = _zz_904[88];
  assign _zz_994 = _zz_904[89];
  assign _zz_995 = _zz_904[90];
  assign _zz_996 = _zz_904[91];
  assign _zz_997 = _zz_904[92];
  assign _zz_998 = _zz_904[93];
  assign _zz_999 = _zz_904[94];
  assign _zz_1000 = _zz_904[95];
  assign _zz_1001 = _zz_904[96];
  assign _zz_1002 = _zz_904[97];
  assign _zz_1003 = _zz_904[98];
  assign _zz_1004 = _zz_904[99];
  assign _zz_1005 = _zz_904[100];
  assign _zz_1006 = _zz_904[101];
  assign _zz_1007 = _zz_904[102];
  assign _zz_1008 = _zz_904[103];
  assign _zz_1009 = _zz_904[104];
  assign _zz_1010 = _zz_904[105];
  assign _zz_1011 = _zz_904[106];
  assign _zz_1012 = _zz_904[107];
  assign _zz_1013 = _zz_904[108];
  assign _zz_1014 = _zz_904[109];
  assign _zz_1015 = _zz_904[110];
  assign _zz_1016 = _zz_904[111];
  assign _zz_1017 = _zz_904[112];
  assign _zz_1018 = _zz_904[113];
  assign _zz_1019 = _zz_904[114];
  assign _zz_1020 = _zz_904[115];
  assign _zz_1021 = _zz_904[116];
  assign _zz_1022 = _zz_904[117];
  assign _zz_1023 = _zz_904[118];
  assign _zz_1024 = _zz_904[119];
  assign _zz_1025 = _zz_904[120];
  assign _zz_1026 = _zz_904[121];
  assign _zz_1027 = _zz_904[122];
  assign _zz_1028 = _zz_904[123];
  assign _zz_1029 = _zz_904[124];
  assign _zz_1030 = _zz_904[125];
  assign _zz_1031 = _zz_904[126];
  assign _zz_1032 = _zz_904[127];
  assign when_DCache_l217_3 = (is_hit && mru_full);
  assign when_DCache_l224_3 = (is_hit && cache_hit_3);
  assign when_DCache_l227_3 = (next_level_rdone && (2'b11 == evict_id_miss));
  assign when_DCache_l232_3 = (next_level_rdone && (2'b11 == evict_id_miss));
  assign when_DCache_l237_3 = ((flush || is_miss) || is_write);
  assign when_DCache_l240_3 = ((flush_done || next_level_rdone) || next_level_wdone);
  assign _zz_cpu_rsp_payload_data = _zz__zz_cpu_rsp_payload_data;
  assign _zz_cpu_rsp_payload_data_1 = _zz__zz_cpu_rsp_payload_data_1;
  assign cpu_rsp_payload_data = (is_hit ? _zz_cpu_rsp_payload_data_2 : _zz_cpu_rsp_payload_data_3);
  assign cpu_rsp_valid = (is_hit ? _zz_cpu_rsp_valid : _zz_cpu_rsp_valid_1);
  assign cpu_cmd_ready = cpu_cmd_ready_1;
  assign stall = (((is_miss || is_write) || (! cpu_cmd_ready_1)) && (! next_level_wdone));
  assign next_level_cmd_payload_addr = (cpu_cmd_payload_wen ? {cpu_cmd_payload_addr[63 : 3],3'b000} : {cpu_cmd_payload_addr[63 : 6],6'h0});
  assign next_level_cmd_payload_len = (cpu_cmd_payload_wen ? 4'b0000 : 4'b0111);
  assign next_level_cmd_payload_size = 3'b011;
  assign next_level_cmd_payload_wen = cpu_cmd_payload_wen;
  assign next_level_cmd_payload_wdata = next_level_wdata;
  assign next_level_cmd_payload_wstrb = next_level_wstrb;
  assign next_level_cmd_valid = next_level_cmd_valid_1;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      ways_0_metas_0_vld <= 1'b0;
      ways_0_metas_0_tag <= 51'h0;
      ways_0_metas_0_mru <= 1'b0;
      ways_0_metas_1_vld <= 1'b0;
      ways_0_metas_1_tag <= 51'h0;
      ways_0_metas_1_mru <= 1'b0;
      ways_0_metas_2_vld <= 1'b0;
      ways_0_metas_2_tag <= 51'h0;
      ways_0_metas_2_mru <= 1'b0;
      ways_0_metas_3_vld <= 1'b0;
      ways_0_metas_3_tag <= 51'h0;
      ways_0_metas_3_mru <= 1'b0;
      ways_0_metas_4_vld <= 1'b0;
      ways_0_metas_4_tag <= 51'h0;
      ways_0_metas_4_mru <= 1'b0;
      ways_0_metas_5_vld <= 1'b0;
      ways_0_metas_5_tag <= 51'h0;
      ways_0_metas_5_mru <= 1'b0;
      ways_0_metas_6_vld <= 1'b0;
      ways_0_metas_6_tag <= 51'h0;
      ways_0_metas_6_mru <= 1'b0;
      ways_0_metas_7_vld <= 1'b0;
      ways_0_metas_7_tag <= 51'h0;
      ways_0_metas_7_mru <= 1'b0;
      ways_0_metas_8_vld <= 1'b0;
      ways_0_metas_8_tag <= 51'h0;
      ways_0_metas_8_mru <= 1'b0;
      ways_0_metas_9_vld <= 1'b0;
      ways_0_metas_9_tag <= 51'h0;
      ways_0_metas_9_mru <= 1'b0;
      ways_0_metas_10_vld <= 1'b0;
      ways_0_metas_10_tag <= 51'h0;
      ways_0_metas_10_mru <= 1'b0;
      ways_0_metas_11_vld <= 1'b0;
      ways_0_metas_11_tag <= 51'h0;
      ways_0_metas_11_mru <= 1'b0;
      ways_0_metas_12_vld <= 1'b0;
      ways_0_metas_12_tag <= 51'h0;
      ways_0_metas_12_mru <= 1'b0;
      ways_0_metas_13_vld <= 1'b0;
      ways_0_metas_13_tag <= 51'h0;
      ways_0_metas_13_mru <= 1'b0;
      ways_0_metas_14_vld <= 1'b0;
      ways_0_metas_14_tag <= 51'h0;
      ways_0_metas_14_mru <= 1'b0;
      ways_0_metas_15_vld <= 1'b0;
      ways_0_metas_15_tag <= 51'h0;
      ways_0_metas_15_mru <= 1'b0;
      ways_0_metas_16_vld <= 1'b0;
      ways_0_metas_16_tag <= 51'h0;
      ways_0_metas_16_mru <= 1'b0;
      ways_0_metas_17_vld <= 1'b0;
      ways_0_metas_17_tag <= 51'h0;
      ways_0_metas_17_mru <= 1'b0;
      ways_0_metas_18_vld <= 1'b0;
      ways_0_metas_18_tag <= 51'h0;
      ways_0_metas_18_mru <= 1'b0;
      ways_0_metas_19_vld <= 1'b0;
      ways_0_metas_19_tag <= 51'h0;
      ways_0_metas_19_mru <= 1'b0;
      ways_0_metas_20_vld <= 1'b0;
      ways_0_metas_20_tag <= 51'h0;
      ways_0_metas_20_mru <= 1'b0;
      ways_0_metas_21_vld <= 1'b0;
      ways_0_metas_21_tag <= 51'h0;
      ways_0_metas_21_mru <= 1'b0;
      ways_0_metas_22_vld <= 1'b0;
      ways_0_metas_22_tag <= 51'h0;
      ways_0_metas_22_mru <= 1'b0;
      ways_0_metas_23_vld <= 1'b0;
      ways_0_metas_23_tag <= 51'h0;
      ways_0_metas_23_mru <= 1'b0;
      ways_0_metas_24_vld <= 1'b0;
      ways_0_metas_24_tag <= 51'h0;
      ways_0_metas_24_mru <= 1'b0;
      ways_0_metas_25_vld <= 1'b0;
      ways_0_metas_25_tag <= 51'h0;
      ways_0_metas_25_mru <= 1'b0;
      ways_0_metas_26_vld <= 1'b0;
      ways_0_metas_26_tag <= 51'h0;
      ways_0_metas_26_mru <= 1'b0;
      ways_0_metas_27_vld <= 1'b0;
      ways_0_metas_27_tag <= 51'h0;
      ways_0_metas_27_mru <= 1'b0;
      ways_0_metas_28_vld <= 1'b0;
      ways_0_metas_28_tag <= 51'h0;
      ways_0_metas_28_mru <= 1'b0;
      ways_0_metas_29_vld <= 1'b0;
      ways_0_metas_29_tag <= 51'h0;
      ways_0_metas_29_mru <= 1'b0;
      ways_0_metas_30_vld <= 1'b0;
      ways_0_metas_30_tag <= 51'h0;
      ways_0_metas_30_mru <= 1'b0;
      ways_0_metas_31_vld <= 1'b0;
      ways_0_metas_31_tag <= 51'h0;
      ways_0_metas_31_mru <= 1'b0;
      ways_0_metas_32_vld <= 1'b0;
      ways_0_metas_32_tag <= 51'h0;
      ways_0_metas_32_mru <= 1'b0;
      ways_0_metas_33_vld <= 1'b0;
      ways_0_metas_33_tag <= 51'h0;
      ways_0_metas_33_mru <= 1'b0;
      ways_0_metas_34_vld <= 1'b0;
      ways_0_metas_34_tag <= 51'h0;
      ways_0_metas_34_mru <= 1'b0;
      ways_0_metas_35_vld <= 1'b0;
      ways_0_metas_35_tag <= 51'h0;
      ways_0_metas_35_mru <= 1'b0;
      ways_0_metas_36_vld <= 1'b0;
      ways_0_metas_36_tag <= 51'h0;
      ways_0_metas_36_mru <= 1'b0;
      ways_0_metas_37_vld <= 1'b0;
      ways_0_metas_37_tag <= 51'h0;
      ways_0_metas_37_mru <= 1'b0;
      ways_0_metas_38_vld <= 1'b0;
      ways_0_metas_38_tag <= 51'h0;
      ways_0_metas_38_mru <= 1'b0;
      ways_0_metas_39_vld <= 1'b0;
      ways_0_metas_39_tag <= 51'h0;
      ways_0_metas_39_mru <= 1'b0;
      ways_0_metas_40_vld <= 1'b0;
      ways_0_metas_40_tag <= 51'h0;
      ways_0_metas_40_mru <= 1'b0;
      ways_0_metas_41_vld <= 1'b0;
      ways_0_metas_41_tag <= 51'h0;
      ways_0_metas_41_mru <= 1'b0;
      ways_0_metas_42_vld <= 1'b0;
      ways_0_metas_42_tag <= 51'h0;
      ways_0_metas_42_mru <= 1'b0;
      ways_0_metas_43_vld <= 1'b0;
      ways_0_metas_43_tag <= 51'h0;
      ways_0_metas_43_mru <= 1'b0;
      ways_0_metas_44_vld <= 1'b0;
      ways_0_metas_44_tag <= 51'h0;
      ways_0_metas_44_mru <= 1'b0;
      ways_0_metas_45_vld <= 1'b0;
      ways_0_metas_45_tag <= 51'h0;
      ways_0_metas_45_mru <= 1'b0;
      ways_0_metas_46_vld <= 1'b0;
      ways_0_metas_46_tag <= 51'h0;
      ways_0_metas_46_mru <= 1'b0;
      ways_0_metas_47_vld <= 1'b0;
      ways_0_metas_47_tag <= 51'h0;
      ways_0_metas_47_mru <= 1'b0;
      ways_0_metas_48_vld <= 1'b0;
      ways_0_metas_48_tag <= 51'h0;
      ways_0_metas_48_mru <= 1'b0;
      ways_0_metas_49_vld <= 1'b0;
      ways_0_metas_49_tag <= 51'h0;
      ways_0_metas_49_mru <= 1'b0;
      ways_0_metas_50_vld <= 1'b0;
      ways_0_metas_50_tag <= 51'h0;
      ways_0_metas_50_mru <= 1'b0;
      ways_0_metas_51_vld <= 1'b0;
      ways_0_metas_51_tag <= 51'h0;
      ways_0_metas_51_mru <= 1'b0;
      ways_0_metas_52_vld <= 1'b0;
      ways_0_metas_52_tag <= 51'h0;
      ways_0_metas_52_mru <= 1'b0;
      ways_0_metas_53_vld <= 1'b0;
      ways_0_metas_53_tag <= 51'h0;
      ways_0_metas_53_mru <= 1'b0;
      ways_0_metas_54_vld <= 1'b0;
      ways_0_metas_54_tag <= 51'h0;
      ways_0_metas_54_mru <= 1'b0;
      ways_0_metas_55_vld <= 1'b0;
      ways_0_metas_55_tag <= 51'h0;
      ways_0_metas_55_mru <= 1'b0;
      ways_0_metas_56_vld <= 1'b0;
      ways_0_metas_56_tag <= 51'h0;
      ways_0_metas_56_mru <= 1'b0;
      ways_0_metas_57_vld <= 1'b0;
      ways_0_metas_57_tag <= 51'h0;
      ways_0_metas_57_mru <= 1'b0;
      ways_0_metas_58_vld <= 1'b0;
      ways_0_metas_58_tag <= 51'h0;
      ways_0_metas_58_mru <= 1'b0;
      ways_0_metas_59_vld <= 1'b0;
      ways_0_metas_59_tag <= 51'h0;
      ways_0_metas_59_mru <= 1'b0;
      ways_0_metas_60_vld <= 1'b0;
      ways_0_metas_60_tag <= 51'h0;
      ways_0_metas_60_mru <= 1'b0;
      ways_0_metas_61_vld <= 1'b0;
      ways_0_metas_61_tag <= 51'h0;
      ways_0_metas_61_mru <= 1'b0;
      ways_0_metas_62_vld <= 1'b0;
      ways_0_metas_62_tag <= 51'h0;
      ways_0_metas_62_mru <= 1'b0;
      ways_0_metas_63_vld <= 1'b0;
      ways_0_metas_63_tag <= 51'h0;
      ways_0_metas_63_mru <= 1'b0;
      ways_0_metas_64_vld <= 1'b0;
      ways_0_metas_64_tag <= 51'h0;
      ways_0_metas_64_mru <= 1'b0;
      ways_0_metas_65_vld <= 1'b0;
      ways_0_metas_65_tag <= 51'h0;
      ways_0_metas_65_mru <= 1'b0;
      ways_0_metas_66_vld <= 1'b0;
      ways_0_metas_66_tag <= 51'h0;
      ways_0_metas_66_mru <= 1'b0;
      ways_0_metas_67_vld <= 1'b0;
      ways_0_metas_67_tag <= 51'h0;
      ways_0_metas_67_mru <= 1'b0;
      ways_0_metas_68_vld <= 1'b0;
      ways_0_metas_68_tag <= 51'h0;
      ways_0_metas_68_mru <= 1'b0;
      ways_0_metas_69_vld <= 1'b0;
      ways_0_metas_69_tag <= 51'h0;
      ways_0_metas_69_mru <= 1'b0;
      ways_0_metas_70_vld <= 1'b0;
      ways_0_metas_70_tag <= 51'h0;
      ways_0_metas_70_mru <= 1'b0;
      ways_0_metas_71_vld <= 1'b0;
      ways_0_metas_71_tag <= 51'h0;
      ways_0_metas_71_mru <= 1'b0;
      ways_0_metas_72_vld <= 1'b0;
      ways_0_metas_72_tag <= 51'h0;
      ways_0_metas_72_mru <= 1'b0;
      ways_0_metas_73_vld <= 1'b0;
      ways_0_metas_73_tag <= 51'h0;
      ways_0_metas_73_mru <= 1'b0;
      ways_0_metas_74_vld <= 1'b0;
      ways_0_metas_74_tag <= 51'h0;
      ways_0_metas_74_mru <= 1'b0;
      ways_0_metas_75_vld <= 1'b0;
      ways_0_metas_75_tag <= 51'h0;
      ways_0_metas_75_mru <= 1'b0;
      ways_0_metas_76_vld <= 1'b0;
      ways_0_metas_76_tag <= 51'h0;
      ways_0_metas_76_mru <= 1'b0;
      ways_0_metas_77_vld <= 1'b0;
      ways_0_metas_77_tag <= 51'h0;
      ways_0_metas_77_mru <= 1'b0;
      ways_0_metas_78_vld <= 1'b0;
      ways_0_metas_78_tag <= 51'h0;
      ways_0_metas_78_mru <= 1'b0;
      ways_0_metas_79_vld <= 1'b0;
      ways_0_metas_79_tag <= 51'h0;
      ways_0_metas_79_mru <= 1'b0;
      ways_0_metas_80_vld <= 1'b0;
      ways_0_metas_80_tag <= 51'h0;
      ways_0_metas_80_mru <= 1'b0;
      ways_0_metas_81_vld <= 1'b0;
      ways_0_metas_81_tag <= 51'h0;
      ways_0_metas_81_mru <= 1'b0;
      ways_0_metas_82_vld <= 1'b0;
      ways_0_metas_82_tag <= 51'h0;
      ways_0_metas_82_mru <= 1'b0;
      ways_0_metas_83_vld <= 1'b0;
      ways_0_metas_83_tag <= 51'h0;
      ways_0_metas_83_mru <= 1'b0;
      ways_0_metas_84_vld <= 1'b0;
      ways_0_metas_84_tag <= 51'h0;
      ways_0_metas_84_mru <= 1'b0;
      ways_0_metas_85_vld <= 1'b0;
      ways_0_metas_85_tag <= 51'h0;
      ways_0_metas_85_mru <= 1'b0;
      ways_0_metas_86_vld <= 1'b0;
      ways_0_metas_86_tag <= 51'h0;
      ways_0_metas_86_mru <= 1'b0;
      ways_0_metas_87_vld <= 1'b0;
      ways_0_metas_87_tag <= 51'h0;
      ways_0_metas_87_mru <= 1'b0;
      ways_0_metas_88_vld <= 1'b0;
      ways_0_metas_88_tag <= 51'h0;
      ways_0_metas_88_mru <= 1'b0;
      ways_0_metas_89_vld <= 1'b0;
      ways_0_metas_89_tag <= 51'h0;
      ways_0_metas_89_mru <= 1'b0;
      ways_0_metas_90_vld <= 1'b0;
      ways_0_metas_90_tag <= 51'h0;
      ways_0_metas_90_mru <= 1'b0;
      ways_0_metas_91_vld <= 1'b0;
      ways_0_metas_91_tag <= 51'h0;
      ways_0_metas_91_mru <= 1'b0;
      ways_0_metas_92_vld <= 1'b0;
      ways_0_metas_92_tag <= 51'h0;
      ways_0_metas_92_mru <= 1'b0;
      ways_0_metas_93_vld <= 1'b0;
      ways_0_metas_93_tag <= 51'h0;
      ways_0_metas_93_mru <= 1'b0;
      ways_0_metas_94_vld <= 1'b0;
      ways_0_metas_94_tag <= 51'h0;
      ways_0_metas_94_mru <= 1'b0;
      ways_0_metas_95_vld <= 1'b0;
      ways_0_metas_95_tag <= 51'h0;
      ways_0_metas_95_mru <= 1'b0;
      ways_0_metas_96_vld <= 1'b0;
      ways_0_metas_96_tag <= 51'h0;
      ways_0_metas_96_mru <= 1'b0;
      ways_0_metas_97_vld <= 1'b0;
      ways_0_metas_97_tag <= 51'h0;
      ways_0_metas_97_mru <= 1'b0;
      ways_0_metas_98_vld <= 1'b0;
      ways_0_metas_98_tag <= 51'h0;
      ways_0_metas_98_mru <= 1'b0;
      ways_0_metas_99_vld <= 1'b0;
      ways_0_metas_99_tag <= 51'h0;
      ways_0_metas_99_mru <= 1'b0;
      ways_0_metas_100_vld <= 1'b0;
      ways_0_metas_100_tag <= 51'h0;
      ways_0_metas_100_mru <= 1'b0;
      ways_0_metas_101_vld <= 1'b0;
      ways_0_metas_101_tag <= 51'h0;
      ways_0_metas_101_mru <= 1'b0;
      ways_0_metas_102_vld <= 1'b0;
      ways_0_metas_102_tag <= 51'h0;
      ways_0_metas_102_mru <= 1'b0;
      ways_0_metas_103_vld <= 1'b0;
      ways_0_metas_103_tag <= 51'h0;
      ways_0_metas_103_mru <= 1'b0;
      ways_0_metas_104_vld <= 1'b0;
      ways_0_metas_104_tag <= 51'h0;
      ways_0_metas_104_mru <= 1'b0;
      ways_0_metas_105_vld <= 1'b0;
      ways_0_metas_105_tag <= 51'h0;
      ways_0_metas_105_mru <= 1'b0;
      ways_0_metas_106_vld <= 1'b0;
      ways_0_metas_106_tag <= 51'h0;
      ways_0_metas_106_mru <= 1'b0;
      ways_0_metas_107_vld <= 1'b0;
      ways_0_metas_107_tag <= 51'h0;
      ways_0_metas_107_mru <= 1'b0;
      ways_0_metas_108_vld <= 1'b0;
      ways_0_metas_108_tag <= 51'h0;
      ways_0_metas_108_mru <= 1'b0;
      ways_0_metas_109_vld <= 1'b0;
      ways_0_metas_109_tag <= 51'h0;
      ways_0_metas_109_mru <= 1'b0;
      ways_0_metas_110_vld <= 1'b0;
      ways_0_metas_110_tag <= 51'h0;
      ways_0_metas_110_mru <= 1'b0;
      ways_0_metas_111_vld <= 1'b0;
      ways_0_metas_111_tag <= 51'h0;
      ways_0_metas_111_mru <= 1'b0;
      ways_0_metas_112_vld <= 1'b0;
      ways_0_metas_112_tag <= 51'h0;
      ways_0_metas_112_mru <= 1'b0;
      ways_0_metas_113_vld <= 1'b0;
      ways_0_metas_113_tag <= 51'h0;
      ways_0_metas_113_mru <= 1'b0;
      ways_0_metas_114_vld <= 1'b0;
      ways_0_metas_114_tag <= 51'h0;
      ways_0_metas_114_mru <= 1'b0;
      ways_0_metas_115_vld <= 1'b0;
      ways_0_metas_115_tag <= 51'h0;
      ways_0_metas_115_mru <= 1'b0;
      ways_0_metas_116_vld <= 1'b0;
      ways_0_metas_116_tag <= 51'h0;
      ways_0_metas_116_mru <= 1'b0;
      ways_0_metas_117_vld <= 1'b0;
      ways_0_metas_117_tag <= 51'h0;
      ways_0_metas_117_mru <= 1'b0;
      ways_0_metas_118_vld <= 1'b0;
      ways_0_metas_118_tag <= 51'h0;
      ways_0_metas_118_mru <= 1'b0;
      ways_0_metas_119_vld <= 1'b0;
      ways_0_metas_119_tag <= 51'h0;
      ways_0_metas_119_mru <= 1'b0;
      ways_0_metas_120_vld <= 1'b0;
      ways_0_metas_120_tag <= 51'h0;
      ways_0_metas_120_mru <= 1'b0;
      ways_0_metas_121_vld <= 1'b0;
      ways_0_metas_121_tag <= 51'h0;
      ways_0_metas_121_mru <= 1'b0;
      ways_0_metas_122_vld <= 1'b0;
      ways_0_metas_122_tag <= 51'h0;
      ways_0_metas_122_mru <= 1'b0;
      ways_0_metas_123_vld <= 1'b0;
      ways_0_metas_123_tag <= 51'h0;
      ways_0_metas_123_mru <= 1'b0;
      ways_0_metas_124_vld <= 1'b0;
      ways_0_metas_124_tag <= 51'h0;
      ways_0_metas_124_mru <= 1'b0;
      ways_0_metas_125_vld <= 1'b0;
      ways_0_metas_125_tag <= 51'h0;
      ways_0_metas_125_mru <= 1'b0;
      ways_0_metas_126_vld <= 1'b0;
      ways_0_metas_126_tag <= 51'h0;
      ways_0_metas_126_mru <= 1'b0;
      ways_0_metas_127_vld <= 1'b0;
      ways_0_metas_127_tag <= 51'h0;
      ways_0_metas_127_mru <= 1'b0;
      ways_1_metas_0_vld <= 1'b0;
      ways_1_metas_0_tag <= 51'h0;
      ways_1_metas_0_mru <= 1'b0;
      ways_1_metas_1_vld <= 1'b0;
      ways_1_metas_1_tag <= 51'h0;
      ways_1_metas_1_mru <= 1'b0;
      ways_1_metas_2_vld <= 1'b0;
      ways_1_metas_2_tag <= 51'h0;
      ways_1_metas_2_mru <= 1'b0;
      ways_1_metas_3_vld <= 1'b0;
      ways_1_metas_3_tag <= 51'h0;
      ways_1_metas_3_mru <= 1'b0;
      ways_1_metas_4_vld <= 1'b0;
      ways_1_metas_4_tag <= 51'h0;
      ways_1_metas_4_mru <= 1'b0;
      ways_1_metas_5_vld <= 1'b0;
      ways_1_metas_5_tag <= 51'h0;
      ways_1_metas_5_mru <= 1'b0;
      ways_1_metas_6_vld <= 1'b0;
      ways_1_metas_6_tag <= 51'h0;
      ways_1_metas_6_mru <= 1'b0;
      ways_1_metas_7_vld <= 1'b0;
      ways_1_metas_7_tag <= 51'h0;
      ways_1_metas_7_mru <= 1'b0;
      ways_1_metas_8_vld <= 1'b0;
      ways_1_metas_8_tag <= 51'h0;
      ways_1_metas_8_mru <= 1'b0;
      ways_1_metas_9_vld <= 1'b0;
      ways_1_metas_9_tag <= 51'h0;
      ways_1_metas_9_mru <= 1'b0;
      ways_1_metas_10_vld <= 1'b0;
      ways_1_metas_10_tag <= 51'h0;
      ways_1_metas_10_mru <= 1'b0;
      ways_1_metas_11_vld <= 1'b0;
      ways_1_metas_11_tag <= 51'h0;
      ways_1_metas_11_mru <= 1'b0;
      ways_1_metas_12_vld <= 1'b0;
      ways_1_metas_12_tag <= 51'h0;
      ways_1_metas_12_mru <= 1'b0;
      ways_1_metas_13_vld <= 1'b0;
      ways_1_metas_13_tag <= 51'h0;
      ways_1_metas_13_mru <= 1'b0;
      ways_1_metas_14_vld <= 1'b0;
      ways_1_metas_14_tag <= 51'h0;
      ways_1_metas_14_mru <= 1'b0;
      ways_1_metas_15_vld <= 1'b0;
      ways_1_metas_15_tag <= 51'h0;
      ways_1_metas_15_mru <= 1'b0;
      ways_1_metas_16_vld <= 1'b0;
      ways_1_metas_16_tag <= 51'h0;
      ways_1_metas_16_mru <= 1'b0;
      ways_1_metas_17_vld <= 1'b0;
      ways_1_metas_17_tag <= 51'h0;
      ways_1_metas_17_mru <= 1'b0;
      ways_1_metas_18_vld <= 1'b0;
      ways_1_metas_18_tag <= 51'h0;
      ways_1_metas_18_mru <= 1'b0;
      ways_1_metas_19_vld <= 1'b0;
      ways_1_metas_19_tag <= 51'h0;
      ways_1_metas_19_mru <= 1'b0;
      ways_1_metas_20_vld <= 1'b0;
      ways_1_metas_20_tag <= 51'h0;
      ways_1_metas_20_mru <= 1'b0;
      ways_1_metas_21_vld <= 1'b0;
      ways_1_metas_21_tag <= 51'h0;
      ways_1_metas_21_mru <= 1'b0;
      ways_1_metas_22_vld <= 1'b0;
      ways_1_metas_22_tag <= 51'h0;
      ways_1_metas_22_mru <= 1'b0;
      ways_1_metas_23_vld <= 1'b0;
      ways_1_metas_23_tag <= 51'h0;
      ways_1_metas_23_mru <= 1'b0;
      ways_1_metas_24_vld <= 1'b0;
      ways_1_metas_24_tag <= 51'h0;
      ways_1_metas_24_mru <= 1'b0;
      ways_1_metas_25_vld <= 1'b0;
      ways_1_metas_25_tag <= 51'h0;
      ways_1_metas_25_mru <= 1'b0;
      ways_1_metas_26_vld <= 1'b0;
      ways_1_metas_26_tag <= 51'h0;
      ways_1_metas_26_mru <= 1'b0;
      ways_1_metas_27_vld <= 1'b0;
      ways_1_metas_27_tag <= 51'h0;
      ways_1_metas_27_mru <= 1'b0;
      ways_1_metas_28_vld <= 1'b0;
      ways_1_metas_28_tag <= 51'h0;
      ways_1_metas_28_mru <= 1'b0;
      ways_1_metas_29_vld <= 1'b0;
      ways_1_metas_29_tag <= 51'h0;
      ways_1_metas_29_mru <= 1'b0;
      ways_1_metas_30_vld <= 1'b0;
      ways_1_metas_30_tag <= 51'h0;
      ways_1_metas_30_mru <= 1'b0;
      ways_1_metas_31_vld <= 1'b0;
      ways_1_metas_31_tag <= 51'h0;
      ways_1_metas_31_mru <= 1'b0;
      ways_1_metas_32_vld <= 1'b0;
      ways_1_metas_32_tag <= 51'h0;
      ways_1_metas_32_mru <= 1'b0;
      ways_1_metas_33_vld <= 1'b0;
      ways_1_metas_33_tag <= 51'h0;
      ways_1_metas_33_mru <= 1'b0;
      ways_1_metas_34_vld <= 1'b0;
      ways_1_metas_34_tag <= 51'h0;
      ways_1_metas_34_mru <= 1'b0;
      ways_1_metas_35_vld <= 1'b0;
      ways_1_metas_35_tag <= 51'h0;
      ways_1_metas_35_mru <= 1'b0;
      ways_1_metas_36_vld <= 1'b0;
      ways_1_metas_36_tag <= 51'h0;
      ways_1_metas_36_mru <= 1'b0;
      ways_1_metas_37_vld <= 1'b0;
      ways_1_metas_37_tag <= 51'h0;
      ways_1_metas_37_mru <= 1'b0;
      ways_1_metas_38_vld <= 1'b0;
      ways_1_metas_38_tag <= 51'h0;
      ways_1_metas_38_mru <= 1'b0;
      ways_1_metas_39_vld <= 1'b0;
      ways_1_metas_39_tag <= 51'h0;
      ways_1_metas_39_mru <= 1'b0;
      ways_1_metas_40_vld <= 1'b0;
      ways_1_metas_40_tag <= 51'h0;
      ways_1_metas_40_mru <= 1'b0;
      ways_1_metas_41_vld <= 1'b0;
      ways_1_metas_41_tag <= 51'h0;
      ways_1_metas_41_mru <= 1'b0;
      ways_1_metas_42_vld <= 1'b0;
      ways_1_metas_42_tag <= 51'h0;
      ways_1_metas_42_mru <= 1'b0;
      ways_1_metas_43_vld <= 1'b0;
      ways_1_metas_43_tag <= 51'h0;
      ways_1_metas_43_mru <= 1'b0;
      ways_1_metas_44_vld <= 1'b0;
      ways_1_metas_44_tag <= 51'h0;
      ways_1_metas_44_mru <= 1'b0;
      ways_1_metas_45_vld <= 1'b0;
      ways_1_metas_45_tag <= 51'h0;
      ways_1_metas_45_mru <= 1'b0;
      ways_1_metas_46_vld <= 1'b0;
      ways_1_metas_46_tag <= 51'h0;
      ways_1_metas_46_mru <= 1'b0;
      ways_1_metas_47_vld <= 1'b0;
      ways_1_metas_47_tag <= 51'h0;
      ways_1_metas_47_mru <= 1'b0;
      ways_1_metas_48_vld <= 1'b0;
      ways_1_metas_48_tag <= 51'h0;
      ways_1_metas_48_mru <= 1'b0;
      ways_1_metas_49_vld <= 1'b0;
      ways_1_metas_49_tag <= 51'h0;
      ways_1_metas_49_mru <= 1'b0;
      ways_1_metas_50_vld <= 1'b0;
      ways_1_metas_50_tag <= 51'h0;
      ways_1_metas_50_mru <= 1'b0;
      ways_1_metas_51_vld <= 1'b0;
      ways_1_metas_51_tag <= 51'h0;
      ways_1_metas_51_mru <= 1'b0;
      ways_1_metas_52_vld <= 1'b0;
      ways_1_metas_52_tag <= 51'h0;
      ways_1_metas_52_mru <= 1'b0;
      ways_1_metas_53_vld <= 1'b0;
      ways_1_metas_53_tag <= 51'h0;
      ways_1_metas_53_mru <= 1'b0;
      ways_1_metas_54_vld <= 1'b0;
      ways_1_metas_54_tag <= 51'h0;
      ways_1_metas_54_mru <= 1'b0;
      ways_1_metas_55_vld <= 1'b0;
      ways_1_metas_55_tag <= 51'h0;
      ways_1_metas_55_mru <= 1'b0;
      ways_1_metas_56_vld <= 1'b0;
      ways_1_metas_56_tag <= 51'h0;
      ways_1_metas_56_mru <= 1'b0;
      ways_1_metas_57_vld <= 1'b0;
      ways_1_metas_57_tag <= 51'h0;
      ways_1_metas_57_mru <= 1'b0;
      ways_1_metas_58_vld <= 1'b0;
      ways_1_metas_58_tag <= 51'h0;
      ways_1_metas_58_mru <= 1'b0;
      ways_1_metas_59_vld <= 1'b0;
      ways_1_metas_59_tag <= 51'h0;
      ways_1_metas_59_mru <= 1'b0;
      ways_1_metas_60_vld <= 1'b0;
      ways_1_metas_60_tag <= 51'h0;
      ways_1_metas_60_mru <= 1'b0;
      ways_1_metas_61_vld <= 1'b0;
      ways_1_metas_61_tag <= 51'h0;
      ways_1_metas_61_mru <= 1'b0;
      ways_1_metas_62_vld <= 1'b0;
      ways_1_metas_62_tag <= 51'h0;
      ways_1_metas_62_mru <= 1'b0;
      ways_1_metas_63_vld <= 1'b0;
      ways_1_metas_63_tag <= 51'h0;
      ways_1_metas_63_mru <= 1'b0;
      ways_1_metas_64_vld <= 1'b0;
      ways_1_metas_64_tag <= 51'h0;
      ways_1_metas_64_mru <= 1'b0;
      ways_1_metas_65_vld <= 1'b0;
      ways_1_metas_65_tag <= 51'h0;
      ways_1_metas_65_mru <= 1'b0;
      ways_1_metas_66_vld <= 1'b0;
      ways_1_metas_66_tag <= 51'h0;
      ways_1_metas_66_mru <= 1'b0;
      ways_1_metas_67_vld <= 1'b0;
      ways_1_metas_67_tag <= 51'h0;
      ways_1_metas_67_mru <= 1'b0;
      ways_1_metas_68_vld <= 1'b0;
      ways_1_metas_68_tag <= 51'h0;
      ways_1_metas_68_mru <= 1'b0;
      ways_1_metas_69_vld <= 1'b0;
      ways_1_metas_69_tag <= 51'h0;
      ways_1_metas_69_mru <= 1'b0;
      ways_1_metas_70_vld <= 1'b0;
      ways_1_metas_70_tag <= 51'h0;
      ways_1_metas_70_mru <= 1'b0;
      ways_1_metas_71_vld <= 1'b0;
      ways_1_metas_71_tag <= 51'h0;
      ways_1_metas_71_mru <= 1'b0;
      ways_1_metas_72_vld <= 1'b0;
      ways_1_metas_72_tag <= 51'h0;
      ways_1_metas_72_mru <= 1'b0;
      ways_1_metas_73_vld <= 1'b0;
      ways_1_metas_73_tag <= 51'h0;
      ways_1_metas_73_mru <= 1'b0;
      ways_1_metas_74_vld <= 1'b0;
      ways_1_metas_74_tag <= 51'h0;
      ways_1_metas_74_mru <= 1'b0;
      ways_1_metas_75_vld <= 1'b0;
      ways_1_metas_75_tag <= 51'h0;
      ways_1_metas_75_mru <= 1'b0;
      ways_1_metas_76_vld <= 1'b0;
      ways_1_metas_76_tag <= 51'h0;
      ways_1_metas_76_mru <= 1'b0;
      ways_1_metas_77_vld <= 1'b0;
      ways_1_metas_77_tag <= 51'h0;
      ways_1_metas_77_mru <= 1'b0;
      ways_1_metas_78_vld <= 1'b0;
      ways_1_metas_78_tag <= 51'h0;
      ways_1_metas_78_mru <= 1'b0;
      ways_1_metas_79_vld <= 1'b0;
      ways_1_metas_79_tag <= 51'h0;
      ways_1_metas_79_mru <= 1'b0;
      ways_1_metas_80_vld <= 1'b0;
      ways_1_metas_80_tag <= 51'h0;
      ways_1_metas_80_mru <= 1'b0;
      ways_1_metas_81_vld <= 1'b0;
      ways_1_metas_81_tag <= 51'h0;
      ways_1_metas_81_mru <= 1'b0;
      ways_1_metas_82_vld <= 1'b0;
      ways_1_metas_82_tag <= 51'h0;
      ways_1_metas_82_mru <= 1'b0;
      ways_1_metas_83_vld <= 1'b0;
      ways_1_metas_83_tag <= 51'h0;
      ways_1_metas_83_mru <= 1'b0;
      ways_1_metas_84_vld <= 1'b0;
      ways_1_metas_84_tag <= 51'h0;
      ways_1_metas_84_mru <= 1'b0;
      ways_1_metas_85_vld <= 1'b0;
      ways_1_metas_85_tag <= 51'h0;
      ways_1_metas_85_mru <= 1'b0;
      ways_1_metas_86_vld <= 1'b0;
      ways_1_metas_86_tag <= 51'h0;
      ways_1_metas_86_mru <= 1'b0;
      ways_1_metas_87_vld <= 1'b0;
      ways_1_metas_87_tag <= 51'h0;
      ways_1_metas_87_mru <= 1'b0;
      ways_1_metas_88_vld <= 1'b0;
      ways_1_metas_88_tag <= 51'h0;
      ways_1_metas_88_mru <= 1'b0;
      ways_1_metas_89_vld <= 1'b0;
      ways_1_metas_89_tag <= 51'h0;
      ways_1_metas_89_mru <= 1'b0;
      ways_1_metas_90_vld <= 1'b0;
      ways_1_metas_90_tag <= 51'h0;
      ways_1_metas_90_mru <= 1'b0;
      ways_1_metas_91_vld <= 1'b0;
      ways_1_metas_91_tag <= 51'h0;
      ways_1_metas_91_mru <= 1'b0;
      ways_1_metas_92_vld <= 1'b0;
      ways_1_metas_92_tag <= 51'h0;
      ways_1_metas_92_mru <= 1'b0;
      ways_1_metas_93_vld <= 1'b0;
      ways_1_metas_93_tag <= 51'h0;
      ways_1_metas_93_mru <= 1'b0;
      ways_1_metas_94_vld <= 1'b0;
      ways_1_metas_94_tag <= 51'h0;
      ways_1_metas_94_mru <= 1'b0;
      ways_1_metas_95_vld <= 1'b0;
      ways_1_metas_95_tag <= 51'h0;
      ways_1_metas_95_mru <= 1'b0;
      ways_1_metas_96_vld <= 1'b0;
      ways_1_metas_96_tag <= 51'h0;
      ways_1_metas_96_mru <= 1'b0;
      ways_1_metas_97_vld <= 1'b0;
      ways_1_metas_97_tag <= 51'h0;
      ways_1_metas_97_mru <= 1'b0;
      ways_1_metas_98_vld <= 1'b0;
      ways_1_metas_98_tag <= 51'h0;
      ways_1_metas_98_mru <= 1'b0;
      ways_1_metas_99_vld <= 1'b0;
      ways_1_metas_99_tag <= 51'h0;
      ways_1_metas_99_mru <= 1'b0;
      ways_1_metas_100_vld <= 1'b0;
      ways_1_metas_100_tag <= 51'h0;
      ways_1_metas_100_mru <= 1'b0;
      ways_1_metas_101_vld <= 1'b0;
      ways_1_metas_101_tag <= 51'h0;
      ways_1_metas_101_mru <= 1'b0;
      ways_1_metas_102_vld <= 1'b0;
      ways_1_metas_102_tag <= 51'h0;
      ways_1_metas_102_mru <= 1'b0;
      ways_1_metas_103_vld <= 1'b0;
      ways_1_metas_103_tag <= 51'h0;
      ways_1_metas_103_mru <= 1'b0;
      ways_1_metas_104_vld <= 1'b0;
      ways_1_metas_104_tag <= 51'h0;
      ways_1_metas_104_mru <= 1'b0;
      ways_1_metas_105_vld <= 1'b0;
      ways_1_metas_105_tag <= 51'h0;
      ways_1_metas_105_mru <= 1'b0;
      ways_1_metas_106_vld <= 1'b0;
      ways_1_metas_106_tag <= 51'h0;
      ways_1_metas_106_mru <= 1'b0;
      ways_1_metas_107_vld <= 1'b0;
      ways_1_metas_107_tag <= 51'h0;
      ways_1_metas_107_mru <= 1'b0;
      ways_1_metas_108_vld <= 1'b0;
      ways_1_metas_108_tag <= 51'h0;
      ways_1_metas_108_mru <= 1'b0;
      ways_1_metas_109_vld <= 1'b0;
      ways_1_metas_109_tag <= 51'h0;
      ways_1_metas_109_mru <= 1'b0;
      ways_1_metas_110_vld <= 1'b0;
      ways_1_metas_110_tag <= 51'h0;
      ways_1_metas_110_mru <= 1'b0;
      ways_1_metas_111_vld <= 1'b0;
      ways_1_metas_111_tag <= 51'h0;
      ways_1_metas_111_mru <= 1'b0;
      ways_1_metas_112_vld <= 1'b0;
      ways_1_metas_112_tag <= 51'h0;
      ways_1_metas_112_mru <= 1'b0;
      ways_1_metas_113_vld <= 1'b0;
      ways_1_metas_113_tag <= 51'h0;
      ways_1_metas_113_mru <= 1'b0;
      ways_1_metas_114_vld <= 1'b0;
      ways_1_metas_114_tag <= 51'h0;
      ways_1_metas_114_mru <= 1'b0;
      ways_1_metas_115_vld <= 1'b0;
      ways_1_metas_115_tag <= 51'h0;
      ways_1_metas_115_mru <= 1'b0;
      ways_1_metas_116_vld <= 1'b0;
      ways_1_metas_116_tag <= 51'h0;
      ways_1_metas_116_mru <= 1'b0;
      ways_1_metas_117_vld <= 1'b0;
      ways_1_metas_117_tag <= 51'h0;
      ways_1_metas_117_mru <= 1'b0;
      ways_1_metas_118_vld <= 1'b0;
      ways_1_metas_118_tag <= 51'h0;
      ways_1_metas_118_mru <= 1'b0;
      ways_1_metas_119_vld <= 1'b0;
      ways_1_metas_119_tag <= 51'h0;
      ways_1_metas_119_mru <= 1'b0;
      ways_1_metas_120_vld <= 1'b0;
      ways_1_metas_120_tag <= 51'h0;
      ways_1_metas_120_mru <= 1'b0;
      ways_1_metas_121_vld <= 1'b0;
      ways_1_metas_121_tag <= 51'h0;
      ways_1_metas_121_mru <= 1'b0;
      ways_1_metas_122_vld <= 1'b0;
      ways_1_metas_122_tag <= 51'h0;
      ways_1_metas_122_mru <= 1'b0;
      ways_1_metas_123_vld <= 1'b0;
      ways_1_metas_123_tag <= 51'h0;
      ways_1_metas_123_mru <= 1'b0;
      ways_1_metas_124_vld <= 1'b0;
      ways_1_metas_124_tag <= 51'h0;
      ways_1_metas_124_mru <= 1'b0;
      ways_1_metas_125_vld <= 1'b0;
      ways_1_metas_125_tag <= 51'h0;
      ways_1_metas_125_mru <= 1'b0;
      ways_1_metas_126_vld <= 1'b0;
      ways_1_metas_126_tag <= 51'h0;
      ways_1_metas_126_mru <= 1'b0;
      ways_1_metas_127_vld <= 1'b0;
      ways_1_metas_127_tag <= 51'h0;
      ways_1_metas_127_mru <= 1'b0;
      ways_2_metas_0_vld <= 1'b0;
      ways_2_metas_0_tag <= 51'h0;
      ways_2_metas_0_mru <= 1'b0;
      ways_2_metas_1_vld <= 1'b0;
      ways_2_metas_1_tag <= 51'h0;
      ways_2_metas_1_mru <= 1'b0;
      ways_2_metas_2_vld <= 1'b0;
      ways_2_metas_2_tag <= 51'h0;
      ways_2_metas_2_mru <= 1'b0;
      ways_2_metas_3_vld <= 1'b0;
      ways_2_metas_3_tag <= 51'h0;
      ways_2_metas_3_mru <= 1'b0;
      ways_2_metas_4_vld <= 1'b0;
      ways_2_metas_4_tag <= 51'h0;
      ways_2_metas_4_mru <= 1'b0;
      ways_2_metas_5_vld <= 1'b0;
      ways_2_metas_5_tag <= 51'h0;
      ways_2_metas_5_mru <= 1'b0;
      ways_2_metas_6_vld <= 1'b0;
      ways_2_metas_6_tag <= 51'h0;
      ways_2_metas_6_mru <= 1'b0;
      ways_2_metas_7_vld <= 1'b0;
      ways_2_metas_7_tag <= 51'h0;
      ways_2_metas_7_mru <= 1'b0;
      ways_2_metas_8_vld <= 1'b0;
      ways_2_metas_8_tag <= 51'h0;
      ways_2_metas_8_mru <= 1'b0;
      ways_2_metas_9_vld <= 1'b0;
      ways_2_metas_9_tag <= 51'h0;
      ways_2_metas_9_mru <= 1'b0;
      ways_2_metas_10_vld <= 1'b0;
      ways_2_metas_10_tag <= 51'h0;
      ways_2_metas_10_mru <= 1'b0;
      ways_2_metas_11_vld <= 1'b0;
      ways_2_metas_11_tag <= 51'h0;
      ways_2_metas_11_mru <= 1'b0;
      ways_2_metas_12_vld <= 1'b0;
      ways_2_metas_12_tag <= 51'h0;
      ways_2_metas_12_mru <= 1'b0;
      ways_2_metas_13_vld <= 1'b0;
      ways_2_metas_13_tag <= 51'h0;
      ways_2_metas_13_mru <= 1'b0;
      ways_2_metas_14_vld <= 1'b0;
      ways_2_metas_14_tag <= 51'h0;
      ways_2_metas_14_mru <= 1'b0;
      ways_2_metas_15_vld <= 1'b0;
      ways_2_metas_15_tag <= 51'h0;
      ways_2_metas_15_mru <= 1'b0;
      ways_2_metas_16_vld <= 1'b0;
      ways_2_metas_16_tag <= 51'h0;
      ways_2_metas_16_mru <= 1'b0;
      ways_2_metas_17_vld <= 1'b0;
      ways_2_metas_17_tag <= 51'h0;
      ways_2_metas_17_mru <= 1'b0;
      ways_2_metas_18_vld <= 1'b0;
      ways_2_metas_18_tag <= 51'h0;
      ways_2_metas_18_mru <= 1'b0;
      ways_2_metas_19_vld <= 1'b0;
      ways_2_metas_19_tag <= 51'h0;
      ways_2_metas_19_mru <= 1'b0;
      ways_2_metas_20_vld <= 1'b0;
      ways_2_metas_20_tag <= 51'h0;
      ways_2_metas_20_mru <= 1'b0;
      ways_2_metas_21_vld <= 1'b0;
      ways_2_metas_21_tag <= 51'h0;
      ways_2_metas_21_mru <= 1'b0;
      ways_2_metas_22_vld <= 1'b0;
      ways_2_metas_22_tag <= 51'h0;
      ways_2_metas_22_mru <= 1'b0;
      ways_2_metas_23_vld <= 1'b0;
      ways_2_metas_23_tag <= 51'h0;
      ways_2_metas_23_mru <= 1'b0;
      ways_2_metas_24_vld <= 1'b0;
      ways_2_metas_24_tag <= 51'h0;
      ways_2_metas_24_mru <= 1'b0;
      ways_2_metas_25_vld <= 1'b0;
      ways_2_metas_25_tag <= 51'h0;
      ways_2_metas_25_mru <= 1'b0;
      ways_2_metas_26_vld <= 1'b0;
      ways_2_metas_26_tag <= 51'h0;
      ways_2_metas_26_mru <= 1'b0;
      ways_2_metas_27_vld <= 1'b0;
      ways_2_metas_27_tag <= 51'h0;
      ways_2_metas_27_mru <= 1'b0;
      ways_2_metas_28_vld <= 1'b0;
      ways_2_metas_28_tag <= 51'h0;
      ways_2_metas_28_mru <= 1'b0;
      ways_2_metas_29_vld <= 1'b0;
      ways_2_metas_29_tag <= 51'h0;
      ways_2_metas_29_mru <= 1'b0;
      ways_2_metas_30_vld <= 1'b0;
      ways_2_metas_30_tag <= 51'h0;
      ways_2_metas_30_mru <= 1'b0;
      ways_2_metas_31_vld <= 1'b0;
      ways_2_metas_31_tag <= 51'h0;
      ways_2_metas_31_mru <= 1'b0;
      ways_2_metas_32_vld <= 1'b0;
      ways_2_metas_32_tag <= 51'h0;
      ways_2_metas_32_mru <= 1'b0;
      ways_2_metas_33_vld <= 1'b0;
      ways_2_metas_33_tag <= 51'h0;
      ways_2_metas_33_mru <= 1'b0;
      ways_2_metas_34_vld <= 1'b0;
      ways_2_metas_34_tag <= 51'h0;
      ways_2_metas_34_mru <= 1'b0;
      ways_2_metas_35_vld <= 1'b0;
      ways_2_metas_35_tag <= 51'h0;
      ways_2_metas_35_mru <= 1'b0;
      ways_2_metas_36_vld <= 1'b0;
      ways_2_metas_36_tag <= 51'h0;
      ways_2_metas_36_mru <= 1'b0;
      ways_2_metas_37_vld <= 1'b0;
      ways_2_metas_37_tag <= 51'h0;
      ways_2_metas_37_mru <= 1'b0;
      ways_2_metas_38_vld <= 1'b0;
      ways_2_metas_38_tag <= 51'h0;
      ways_2_metas_38_mru <= 1'b0;
      ways_2_metas_39_vld <= 1'b0;
      ways_2_metas_39_tag <= 51'h0;
      ways_2_metas_39_mru <= 1'b0;
      ways_2_metas_40_vld <= 1'b0;
      ways_2_metas_40_tag <= 51'h0;
      ways_2_metas_40_mru <= 1'b0;
      ways_2_metas_41_vld <= 1'b0;
      ways_2_metas_41_tag <= 51'h0;
      ways_2_metas_41_mru <= 1'b0;
      ways_2_metas_42_vld <= 1'b0;
      ways_2_metas_42_tag <= 51'h0;
      ways_2_metas_42_mru <= 1'b0;
      ways_2_metas_43_vld <= 1'b0;
      ways_2_metas_43_tag <= 51'h0;
      ways_2_metas_43_mru <= 1'b0;
      ways_2_metas_44_vld <= 1'b0;
      ways_2_metas_44_tag <= 51'h0;
      ways_2_metas_44_mru <= 1'b0;
      ways_2_metas_45_vld <= 1'b0;
      ways_2_metas_45_tag <= 51'h0;
      ways_2_metas_45_mru <= 1'b0;
      ways_2_metas_46_vld <= 1'b0;
      ways_2_metas_46_tag <= 51'h0;
      ways_2_metas_46_mru <= 1'b0;
      ways_2_metas_47_vld <= 1'b0;
      ways_2_metas_47_tag <= 51'h0;
      ways_2_metas_47_mru <= 1'b0;
      ways_2_metas_48_vld <= 1'b0;
      ways_2_metas_48_tag <= 51'h0;
      ways_2_metas_48_mru <= 1'b0;
      ways_2_metas_49_vld <= 1'b0;
      ways_2_metas_49_tag <= 51'h0;
      ways_2_metas_49_mru <= 1'b0;
      ways_2_metas_50_vld <= 1'b0;
      ways_2_metas_50_tag <= 51'h0;
      ways_2_metas_50_mru <= 1'b0;
      ways_2_metas_51_vld <= 1'b0;
      ways_2_metas_51_tag <= 51'h0;
      ways_2_metas_51_mru <= 1'b0;
      ways_2_metas_52_vld <= 1'b0;
      ways_2_metas_52_tag <= 51'h0;
      ways_2_metas_52_mru <= 1'b0;
      ways_2_metas_53_vld <= 1'b0;
      ways_2_metas_53_tag <= 51'h0;
      ways_2_metas_53_mru <= 1'b0;
      ways_2_metas_54_vld <= 1'b0;
      ways_2_metas_54_tag <= 51'h0;
      ways_2_metas_54_mru <= 1'b0;
      ways_2_metas_55_vld <= 1'b0;
      ways_2_metas_55_tag <= 51'h0;
      ways_2_metas_55_mru <= 1'b0;
      ways_2_metas_56_vld <= 1'b0;
      ways_2_metas_56_tag <= 51'h0;
      ways_2_metas_56_mru <= 1'b0;
      ways_2_metas_57_vld <= 1'b0;
      ways_2_metas_57_tag <= 51'h0;
      ways_2_metas_57_mru <= 1'b0;
      ways_2_metas_58_vld <= 1'b0;
      ways_2_metas_58_tag <= 51'h0;
      ways_2_metas_58_mru <= 1'b0;
      ways_2_metas_59_vld <= 1'b0;
      ways_2_metas_59_tag <= 51'h0;
      ways_2_metas_59_mru <= 1'b0;
      ways_2_metas_60_vld <= 1'b0;
      ways_2_metas_60_tag <= 51'h0;
      ways_2_metas_60_mru <= 1'b0;
      ways_2_metas_61_vld <= 1'b0;
      ways_2_metas_61_tag <= 51'h0;
      ways_2_metas_61_mru <= 1'b0;
      ways_2_metas_62_vld <= 1'b0;
      ways_2_metas_62_tag <= 51'h0;
      ways_2_metas_62_mru <= 1'b0;
      ways_2_metas_63_vld <= 1'b0;
      ways_2_metas_63_tag <= 51'h0;
      ways_2_metas_63_mru <= 1'b0;
      ways_2_metas_64_vld <= 1'b0;
      ways_2_metas_64_tag <= 51'h0;
      ways_2_metas_64_mru <= 1'b0;
      ways_2_metas_65_vld <= 1'b0;
      ways_2_metas_65_tag <= 51'h0;
      ways_2_metas_65_mru <= 1'b0;
      ways_2_metas_66_vld <= 1'b0;
      ways_2_metas_66_tag <= 51'h0;
      ways_2_metas_66_mru <= 1'b0;
      ways_2_metas_67_vld <= 1'b0;
      ways_2_metas_67_tag <= 51'h0;
      ways_2_metas_67_mru <= 1'b0;
      ways_2_metas_68_vld <= 1'b0;
      ways_2_metas_68_tag <= 51'h0;
      ways_2_metas_68_mru <= 1'b0;
      ways_2_metas_69_vld <= 1'b0;
      ways_2_metas_69_tag <= 51'h0;
      ways_2_metas_69_mru <= 1'b0;
      ways_2_metas_70_vld <= 1'b0;
      ways_2_metas_70_tag <= 51'h0;
      ways_2_metas_70_mru <= 1'b0;
      ways_2_metas_71_vld <= 1'b0;
      ways_2_metas_71_tag <= 51'h0;
      ways_2_metas_71_mru <= 1'b0;
      ways_2_metas_72_vld <= 1'b0;
      ways_2_metas_72_tag <= 51'h0;
      ways_2_metas_72_mru <= 1'b0;
      ways_2_metas_73_vld <= 1'b0;
      ways_2_metas_73_tag <= 51'h0;
      ways_2_metas_73_mru <= 1'b0;
      ways_2_metas_74_vld <= 1'b0;
      ways_2_metas_74_tag <= 51'h0;
      ways_2_metas_74_mru <= 1'b0;
      ways_2_metas_75_vld <= 1'b0;
      ways_2_metas_75_tag <= 51'h0;
      ways_2_metas_75_mru <= 1'b0;
      ways_2_metas_76_vld <= 1'b0;
      ways_2_metas_76_tag <= 51'h0;
      ways_2_metas_76_mru <= 1'b0;
      ways_2_metas_77_vld <= 1'b0;
      ways_2_metas_77_tag <= 51'h0;
      ways_2_metas_77_mru <= 1'b0;
      ways_2_metas_78_vld <= 1'b0;
      ways_2_metas_78_tag <= 51'h0;
      ways_2_metas_78_mru <= 1'b0;
      ways_2_metas_79_vld <= 1'b0;
      ways_2_metas_79_tag <= 51'h0;
      ways_2_metas_79_mru <= 1'b0;
      ways_2_metas_80_vld <= 1'b0;
      ways_2_metas_80_tag <= 51'h0;
      ways_2_metas_80_mru <= 1'b0;
      ways_2_metas_81_vld <= 1'b0;
      ways_2_metas_81_tag <= 51'h0;
      ways_2_metas_81_mru <= 1'b0;
      ways_2_metas_82_vld <= 1'b0;
      ways_2_metas_82_tag <= 51'h0;
      ways_2_metas_82_mru <= 1'b0;
      ways_2_metas_83_vld <= 1'b0;
      ways_2_metas_83_tag <= 51'h0;
      ways_2_metas_83_mru <= 1'b0;
      ways_2_metas_84_vld <= 1'b0;
      ways_2_metas_84_tag <= 51'h0;
      ways_2_metas_84_mru <= 1'b0;
      ways_2_metas_85_vld <= 1'b0;
      ways_2_metas_85_tag <= 51'h0;
      ways_2_metas_85_mru <= 1'b0;
      ways_2_metas_86_vld <= 1'b0;
      ways_2_metas_86_tag <= 51'h0;
      ways_2_metas_86_mru <= 1'b0;
      ways_2_metas_87_vld <= 1'b0;
      ways_2_metas_87_tag <= 51'h0;
      ways_2_metas_87_mru <= 1'b0;
      ways_2_metas_88_vld <= 1'b0;
      ways_2_metas_88_tag <= 51'h0;
      ways_2_metas_88_mru <= 1'b0;
      ways_2_metas_89_vld <= 1'b0;
      ways_2_metas_89_tag <= 51'h0;
      ways_2_metas_89_mru <= 1'b0;
      ways_2_metas_90_vld <= 1'b0;
      ways_2_metas_90_tag <= 51'h0;
      ways_2_metas_90_mru <= 1'b0;
      ways_2_metas_91_vld <= 1'b0;
      ways_2_metas_91_tag <= 51'h0;
      ways_2_metas_91_mru <= 1'b0;
      ways_2_metas_92_vld <= 1'b0;
      ways_2_metas_92_tag <= 51'h0;
      ways_2_metas_92_mru <= 1'b0;
      ways_2_metas_93_vld <= 1'b0;
      ways_2_metas_93_tag <= 51'h0;
      ways_2_metas_93_mru <= 1'b0;
      ways_2_metas_94_vld <= 1'b0;
      ways_2_metas_94_tag <= 51'h0;
      ways_2_metas_94_mru <= 1'b0;
      ways_2_metas_95_vld <= 1'b0;
      ways_2_metas_95_tag <= 51'h0;
      ways_2_metas_95_mru <= 1'b0;
      ways_2_metas_96_vld <= 1'b0;
      ways_2_metas_96_tag <= 51'h0;
      ways_2_metas_96_mru <= 1'b0;
      ways_2_metas_97_vld <= 1'b0;
      ways_2_metas_97_tag <= 51'h0;
      ways_2_metas_97_mru <= 1'b0;
      ways_2_metas_98_vld <= 1'b0;
      ways_2_metas_98_tag <= 51'h0;
      ways_2_metas_98_mru <= 1'b0;
      ways_2_metas_99_vld <= 1'b0;
      ways_2_metas_99_tag <= 51'h0;
      ways_2_metas_99_mru <= 1'b0;
      ways_2_metas_100_vld <= 1'b0;
      ways_2_metas_100_tag <= 51'h0;
      ways_2_metas_100_mru <= 1'b0;
      ways_2_metas_101_vld <= 1'b0;
      ways_2_metas_101_tag <= 51'h0;
      ways_2_metas_101_mru <= 1'b0;
      ways_2_metas_102_vld <= 1'b0;
      ways_2_metas_102_tag <= 51'h0;
      ways_2_metas_102_mru <= 1'b0;
      ways_2_metas_103_vld <= 1'b0;
      ways_2_metas_103_tag <= 51'h0;
      ways_2_metas_103_mru <= 1'b0;
      ways_2_metas_104_vld <= 1'b0;
      ways_2_metas_104_tag <= 51'h0;
      ways_2_metas_104_mru <= 1'b0;
      ways_2_metas_105_vld <= 1'b0;
      ways_2_metas_105_tag <= 51'h0;
      ways_2_metas_105_mru <= 1'b0;
      ways_2_metas_106_vld <= 1'b0;
      ways_2_metas_106_tag <= 51'h0;
      ways_2_metas_106_mru <= 1'b0;
      ways_2_metas_107_vld <= 1'b0;
      ways_2_metas_107_tag <= 51'h0;
      ways_2_metas_107_mru <= 1'b0;
      ways_2_metas_108_vld <= 1'b0;
      ways_2_metas_108_tag <= 51'h0;
      ways_2_metas_108_mru <= 1'b0;
      ways_2_metas_109_vld <= 1'b0;
      ways_2_metas_109_tag <= 51'h0;
      ways_2_metas_109_mru <= 1'b0;
      ways_2_metas_110_vld <= 1'b0;
      ways_2_metas_110_tag <= 51'h0;
      ways_2_metas_110_mru <= 1'b0;
      ways_2_metas_111_vld <= 1'b0;
      ways_2_metas_111_tag <= 51'h0;
      ways_2_metas_111_mru <= 1'b0;
      ways_2_metas_112_vld <= 1'b0;
      ways_2_metas_112_tag <= 51'h0;
      ways_2_metas_112_mru <= 1'b0;
      ways_2_metas_113_vld <= 1'b0;
      ways_2_metas_113_tag <= 51'h0;
      ways_2_metas_113_mru <= 1'b0;
      ways_2_metas_114_vld <= 1'b0;
      ways_2_metas_114_tag <= 51'h0;
      ways_2_metas_114_mru <= 1'b0;
      ways_2_metas_115_vld <= 1'b0;
      ways_2_metas_115_tag <= 51'h0;
      ways_2_metas_115_mru <= 1'b0;
      ways_2_metas_116_vld <= 1'b0;
      ways_2_metas_116_tag <= 51'h0;
      ways_2_metas_116_mru <= 1'b0;
      ways_2_metas_117_vld <= 1'b0;
      ways_2_metas_117_tag <= 51'h0;
      ways_2_metas_117_mru <= 1'b0;
      ways_2_metas_118_vld <= 1'b0;
      ways_2_metas_118_tag <= 51'h0;
      ways_2_metas_118_mru <= 1'b0;
      ways_2_metas_119_vld <= 1'b0;
      ways_2_metas_119_tag <= 51'h0;
      ways_2_metas_119_mru <= 1'b0;
      ways_2_metas_120_vld <= 1'b0;
      ways_2_metas_120_tag <= 51'h0;
      ways_2_metas_120_mru <= 1'b0;
      ways_2_metas_121_vld <= 1'b0;
      ways_2_metas_121_tag <= 51'h0;
      ways_2_metas_121_mru <= 1'b0;
      ways_2_metas_122_vld <= 1'b0;
      ways_2_metas_122_tag <= 51'h0;
      ways_2_metas_122_mru <= 1'b0;
      ways_2_metas_123_vld <= 1'b0;
      ways_2_metas_123_tag <= 51'h0;
      ways_2_metas_123_mru <= 1'b0;
      ways_2_metas_124_vld <= 1'b0;
      ways_2_metas_124_tag <= 51'h0;
      ways_2_metas_124_mru <= 1'b0;
      ways_2_metas_125_vld <= 1'b0;
      ways_2_metas_125_tag <= 51'h0;
      ways_2_metas_125_mru <= 1'b0;
      ways_2_metas_126_vld <= 1'b0;
      ways_2_metas_126_tag <= 51'h0;
      ways_2_metas_126_mru <= 1'b0;
      ways_2_metas_127_vld <= 1'b0;
      ways_2_metas_127_tag <= 51'h0;
      ways_2_metas_127_mru <= 1'b0;
      ways_3_metas_0_vld <= 1'b0;
      ways_3_metas_0_tag <= 51'h0;
      ways_3_metas_0_mru <= 1'b0;
      ways_3_metas_1_vld <= 1'b0;
      ways_3_metas_1_tag <= 51'h0;
      ways_3_metas_1_mru <= 1'b0;
      ways_3_metas_2_vld <= 1'b0;
      ways_3_metas_2_tag <= 51'h0;
      ways_3_metas_2_mru <= 1'b0;
      ways_3_metas_3_vld <= 1'b0;
      ways_3_metas_3_tag <= 51'h0;
      ways_3_metas_3_mru <= 1'b0;
      ways_3_metas_4_vld <= 1'b0;
      ways_3_metas_4_tag <= 51'h0;
      ways_3_metas_4_mru <= 1'b0;
      ways_3_metas_5_vld <= 1'b0;
      ways_3_metas_5_tag <= 51'h0;
      ways_3_metas_5_mru <= 1'b0;
      ways_3_metas_6_vld <= 1'b0;
      ways_3_metas_6_tag <= 51'h0;
      ways_3_metas_6_mru <= 1'b0;
      ways_3_metas_7_vld <= 1'b0;
      ways_3_metas_7_tag <= 51'h0;
      ways_3_metas_7_mru <= 1'b0;
      ways_3_metas_8_vld <= 1'b0;
      ways_3_metas_8_tag <= 51'h0;
      ways_3_metas_8_mru <= 1'b0;
      ways_3_metas_9_vld <= 1'b0;
      ways_3_metas_9_tag <= 51'h0;
      ways_3_metas_9_mru <= 1'b0;
      ways_3_metas_10_vld <= 1'b0;
      ways_3_metas_10_tag <= 51'h0;
      ways_3_metas_10_mru <= 1'b0;
      ways_3_metas_11_vld <= 1'b0;
      ways_3_metas_11_tag <= 51'h0;
      ways_3_metas_11_mru <= 1'b0;
      ways_3_metas_12_vld <= 1'b0;
      ways_3_metas_12_tag <= 51'h0;
      ways_3_metas_12_mru <= 1'b0;
      ways_3_metas_13_vld <= 1'b0;
      ways_3_metas_13_tag <= 51'h0;
      ways_3_metas_13_mru <= 1'b0;
      ways_3_metas_14_vld <= 1'b0;
      ways_3_metas_14_tag <= 51'h0;
      ways_3_metas_14_mru <= 1'b0;
      ways_3_metas_15_vld <= 1'b0;
      ways_3_metas_15_tag <= 51'h0;
      ways_3_metas_15_mru <= 1'b0;
      ways_3_metas_16_vld <= 1'b0;
      ways_3_metas_16_tag <= 51'h0;
      ways_3_metas_16_mru <= 1'b0;
      ways_3_metas_17_vld <= 1'b0;
      ways_3_metas_17_tag <= 51'h0;
      ways_3_metas_17_mru <= 1'b0;
      ways_3_metas_18_vld <= 1'b0;
      ways_3_metas_18_tag <= 51'h0;
      ways_3_metas_18_mru <= 1'b0;
      ways_3_metas_19_vld <= 1'b0;
      ways_3_metas_19_tag <= 51'h0;
      ways_3_metas_19_mru <= 1'b0;
      ways_3_metas_20_vld <= 1'b0;
      ways_3_metas_20_tag <= 51'h0;
      ways_3_metas_20_mru <= 1'b0;
      ways_3_metas_21_vld <= 1'b0;
      ways_3_metas_21_tag <= 51'h0;
      ways_3_metas_21_mru <= 1'b0;
      ways_3_metas_22_vld <= 1'b0;
      ways_3_metas_22_tag <= 51'h0;
      ways_3_metas_22_mru <= 1'b0;
      ways_3_metas_23_vld <= 1'b0;
      ways_3_metas_23_tag <= 51'h0;
      ways_3_metas_23_mru <= 1'b0;
      ways_3_metas_24_vld <= 1'b0;
      ways_3_metas_24_tag <= 51'h0;
      ways_3_metas_24_mru <= 1'b0;
      ways_3_metas_25_vld <= 1'b0;
      ways_3_metas_25_tag <= 51'h0;
      ways_3_metas_25_mru <= 1'b0;
      ways_3_metas_26_vld <= 1'b0;
      ways_3_metas_26_tag <= 51'h0;
      ways_3_metas_26_mru <= 1'b0;
      ways_3_metas_27_vld <= 1'b0;
      ways_3_metas_27_tag <= 51'h0;
      ways_3_metas_27_mru <= 1'b0;
      ways_3_metas_28_vld <= 1'b0;
      ways_3_metas_28_tag <= 51'h0;
      ways_3_metas_28_mru <= 1'b0;
      ways_3_metas_29_vld <= 1'b0;
      ways_3_metas_29_tag <= 51'h0;
      ways_3_metas_29_mru <= 1'b0;
      ways_3_metas_30_vld <= 1'b0;
      ways_3_metas_30_tag <= 51'h0;
      ways_3_metas_30_mru <= 1'b0;
      ways_3_metas_31_vld <= 1'b0;
      ways_3_metas_31_tag <= 51'h0;
      ways_3_metas_31_mru <= 1'b0;
      ways_3_metas_32_vld <= 1'b0;
      ways_3_metas_32_tag <= 51'h0;
      ways_3_metas_32_mru <= 1'b0;
      ways_3_metas_33_vld <= 1'b0;
      ways_3_metas_33_tag <= 51'h0;
      ways_3_metas_33_mru <= 1'b0;
      ways_3_metas_34_vld <= 1'b0;
      ways_3_metas_34_tag <= 51'h0;
      ways_3_metas_34_mru <= 1'b0;
      ways_3_metas_35_vld <= 1'b0;
      ways_3_metas_35_tag <= 51'h0;
      ways_3_metas_35_mru <= 1'b0;
      ways_3_metas_36_vld <= 1'b0;
      ways_3_metas_36_tag <= 51'h0;
      ways_3_metas_36_mru <= 1'b0;
      ways_3_metas_37_vld <= 1'b0;
      ways_3_metas_37_tag <= 51'h0;
      ways_3_metas_37_mru <= 1'b0;
      ways_3_metas_38_vld <= 1'b0;
      ways_3_metas_38_tag <= 51'h0;
      ways_3_metas_38_mru <= 1'b0;
      ways_3_metas_39_vld <= 1'b0;
      ways_3_metas_39_tag <= 51'h0;
      ways_3_metas_39_mru <= 1'b0;
      ways_3_metas_40_vld <= 1'b0;
      ways_3_metas_40_tag <= 51'h0;
      ways_3_metas_40_mru <= 1'b0;
      ways_3_metas_41_vld <= 1'b0;
      ways_3_metas_41_tag <= 51'h0;
      ways_3_metas_41_mru <= 1'b0;
      ways_3_metas_42_vld <= 1'b0;
      ways_3_metas_42_tag <= 51'h0;
      ways_3_metas_42_mru <= 1'b0;
      ways_3_metas_43_vld <= 1'b0;
      ways_3_metas_43_tag <= 51'h0;
      ways_3_metas_43_mru <= 1'b0;
      ways_3_metas_44_vld <= 1'b0;
      ways_3_metas_44_tag <= 51'h0;
      ways_3_metas_44_mru <= 1'b0;
      ways_3_metas_45_vld <= 1'b0;
      ways_3_metas_45_tag <= 51'h0;
      ways_3_metas_45_mru <= 1'b0;
      ways_3_metas_46_vld <= 1'b0;
      ways_3_metas_46_tag <= 51'h0;
      ways_3_metas_46_mru <= 1'b0;
      ways_3_metas_47_vld <= 1'b0;
      ways_3_metas_47_tag <= 51'h0;
      ways_3_metas_47_mru <= 1'b0;
      ways_3_metas_48_vld <= 1'b0;
      ways_3_metas_48_tag <= 51'h0;
      ways_3_metas_48_mru <= 1'b0;
      ways_3_metas_49_vld <= 1'b0;
      ways_3_metas_49_tag <= 51'h0;
      ways_3_metas_49_mru <= 1'b0;
      ways_3_metas_50_vld <= 1'b0;
      ways_3_metas_50_tag <= 51'h0;
      ways_3_metas_50_mru <= 1'b0;
      ways_3_metas_51_vld <= 1'b0;
      ways_3_metas_51_tag <= 51'h0;
      ways_3_metas_51_mru <= 1'b0;
      ways_3_metas_52_vld <= 1'b0;
      ways_3_metas_52_tag <= 51'h0;
      ways_3_metas_52_mru <= 1'b0;
      ways_3_metas_53_vld <= 1'b0;
      ways_3_metas_53_tag <= 51'h0;
      ways_3_metas_53_mru <= 1'b0;
      ways_3_metas_54_vld <= 1'b0;
      ways_3_metas_54_tag <= 51'h0;
      ways_3_metas_54_mru <= 1'b0;
      ways_3_metas_55_vld <= 1'b0;
      ways_3_metas_55_tag <= 51'h0;
      ways_3_metas_55_mru <= 1'b0;
      ways_3_metas_56_vld <= 1'b0;
      ways_3_metas_56_tag <= 51'h0;
      ways_3_metas_56_mru <= 1'b0;
      ways_3_metas_57_vld <= 1'b0;
      ways_3_metas_57_tag <= 51'h0;
      ways_3_metas_57_mru <= 1'b0;
      ways_3_metas_58_vld <= 1'b0;
      ways_3_metas_58_tag <= 51'h0;
      ways_3_metas_58_mru <= 1'b0;
      ways_3_metas_59_vld <= 1'b0;
      ways_3_metas_59_tag <= 51'h0;
      ways_3_metas_59_mru <= 1'b0;
      ways_3_metas_60_vld <= 1'b0;
      ways_3_metas_60_tag <= 51'h0;
      ways_3_metas_60_mru <= 1'b0;
      ways_3_metas_61_vld <= 1'b0;
      ways_3_metas_61_tag <= 51'h0;
      ways_3_metas_61_mru <= 1'b0;
      ways_3_metas_62_vld <= 1'b0;
      ways_3_metas_62_tag <= 51'h0;
      ways_3_metas_62_mru <= 1'b0;
      ways_3_metas_63_vld <= 1'b0;
      ways_3_metas_63_tag <= 51'h0;
      ways_3_metas_63_mru <= 1'b0;
      ways_3_metas_64_vld <= 1'b0;
      ways_3_metas_64_tag <= 51'h0;
      ways_3_metas_64_mru <= 1'b0;
      ways_3_metas_65_vld <= 1'b0;
      ways_3_metas_65_tag <= 51'h0;
      ways_3_metas_65_mru <= 1'b0;
      ways_3_metas_66_vld <= 1'b0;
      ways_3_metas_66_tag <= 51'h0;
      ways_3_metas_66_mru <= 1'b0;
      ways_3_metas_67_vld <= 1'b0;
      ways_3_metas_67_tag <= 51'h0;
      ways_3_metas_67_mru <= 1'b0;
      ways_3_metas_68_vld <= 1'b0;
      ways_3_metas_68_tag <= 51'h0;
      ways_3_metas_68_mru <= 1'b0;
      ways_3_metas_69_vld <= 1'b0;
      ways_3_metas_69_tag <= 51'h0;
      ways_3_metas_69_mru <= 1'b0;
      ways_3_metas_70_vld <= 1'b0;
      ways_3_metas_70_tag <= 51'h0;
      ways_3_metas_70_mru <= 1'b0;
      ways_3_metas_71_vld <= 1'b0;
      ways_3_metas_71_tag <= 51'h0;
      ways_3_metas_71_mru <= 1'b0;
      ways_3_metas_72_vld <= 1'b0;
      ways_3_metas_72_tag <= 51'h0;
      ways_3_metas_72_mru <= 1'b0;
      ways_3_metas_73_vld <= 1'b0;
      ways_3_metas_73_tag <= 51'h0;
      ways_3_metas_73_mru <= 1'b0;
      ways_3_metas_74_vld <= 1'b0;
      ways_3_metas_74_tag <= 51'h0;
      ways_3_metas_74_mru <= 1'b0;
      ways_3_metas_75_vld <= 1'b0;
      ways_3_metas_75_tag <= 51'h0;
      ways_3_metas_75_mru <= 1'b0;
      ways_3_metas_76_vld <= 1'b0;
      ways_3_metas_76_tag <= 51'h0;
      ways_3_metas_76_mru <= 1'b0;
      ways_3_metas_77_vld <= 1'b0;
      ways_3_metas_77_tag <= 51'h0;
      ways_3_metas_77_mru <= 1'b0;
      ways_3_metas_78_vld <= 1'b0;
      ways_3_metas_78_tag <= 51'h0;
      ways_3_metas_78_mru <= 1'b0;
      ways_3_metas_79_vld <= 1'b0;
      ways_3_metas_79_tag <= 51'h0;
      ways_3_metas_79_mru <= 1'b0;
      ways_3_metas_80_vld <= 1'b0;
      ways_3_metas_80_tag <= 51'h0;
      ways_3_metas_80_mru <= 1'b0;
      ways_3_metas_81_vld <= 1'b0;
      ways_3_metas_81_tag <= 51'h0;
      ways_3_metas_81_mru <= 1'b0;
      ways_3_metas_82_vld <= 1'b0;
      ways_3_metas_82_tag <= 51'h0;
      ways_3_metas_82_mru <= 1'b0;
      ways_3_metas_83_vld <= 1'b0;
      ways_3_metas_83_tag <= 51'h0;
      ways_3_metas_83_mru <= 1'b0;
      ways_3_metas_84_vld <= 1'b0;
      ways_3_metas_84_tag <= 51'h0;
      ways_3_metas_84_mru <= 1'b0;
      ways_3_metas_85_vld <= 1'b0;
      ways_3_metas_85_tag <= 51'h0;
      ways_3_metas_85_mru <= 1'b0;
      ways_3_metas_86_vld <= 1'b0;
      ways_3_metas_86_tag <= 51'h0;
      ways_3_metas_86_mru <= 1'b0;
      ways_3_metas_87_vld <= 1'b0;
      ways_3_metas_87_tag <= 51'h0;
      ways_3_metas_87_mru <= 1'b0;
      ways_3_metas_88_vld <= 1'b0;
      ways_3_metas_88_tag <= 51'h0;
      ways_3_metas_88_mru <= 1'b0;
      ways_3_metas_89_vld <= 1'b0;
      ways_3_metas_89_tag <= 51'h0;
      ways_3_metas_89_mru <= 1'b0;
      ways_3_metas_90_vld <= 1'b0;
      ways_3_metas_90_tag <= 51'h0;
      ways_3_metas_90_mru <= 1'b0;
      ways_3_metas_91_vld <= 1'b0;
      ways_3_metas_91_tag <= 51'h0;
      ways_3_metas_91_mru <= 1'b0;
      ways_3_metas_92_vld <= 1'b0;
      ways_3_metas_92_tag <= 51'h0;
      ways_3_metas_92_mru <= 1'b0;
      ways_3_metas_93_vld <= 1'b0;
      ways_3_metas_93_tag <= 51'h0;
      ways_3_metas_93_mru <= 1'b0;
      ways_3_metas_94_vld <= 1'b0;
      ways_3_metas_94_tag <= 51'h0;
      ways_3_metas_94_mru <= 1'b0;
      ways_3_metas_95_vld <= 1'b0;
      ways_3_metas_95_tag <= 51'h0;
      ways_3_metas_95_mru <= 1'b0;
      ways_3_metas_96_vld <= 1'b0;
      ways_3_metas_96_tag <= 51'h0;
      ways_3_metas_96_mru <= 1'b0;
      ways_3_metas_97_vld <= 1'b0;
      ways_3_metas_97_tag <= 51'h0;
      ways_3_metas_97_mru <= 1'b0;
      ways_3_metas_98_vld <= 1'b0;
      ways_3_metas_98_tag <= 51'h0;
      ways_3_metas_98_mru <= 1'b0;
      ways_3_metas_99_vld <= 1'b0;
      ways_3_metas_99_tag <= 51'h0;
      ways_3_metas_99_mru <= 1'b0;
      ways_3_metas_100_vld <= 1'b0;
      ways_3_metas_100_tag <= 51'h0;
      ways_3_metas_100_mru <= 1'b0;
      ways_3_metas_101_vld <= 1'b0;
      ways_3_metas_101_tag <= 51'h0;
      ways_3_metas_101_mru <= 1'b0;
      ways_3_metas_102_vld <= 1'b0;
      ways_3_metas_102_tag <= 51'h0;
      ways_3_metas_102_mru <= 1'b0;
      ways_3_metas_103_vld <= 1'b0;
      ways_3_metas_103_tag <= 51'h0;
      ways_3_metas_103_mru <= 1'b0;
      ways_3_metas_104_vld <= 1'b0;
      ways_3_metas_104_tag <= 51'h0;
      ways_3_metas_104_mru <= 1'b0;
      ways_3_metas_105_vld <= 1'b0;
      ways_3_metas_105_tag <= 51'h0;
      ways_3_metas_105_mru <= 1'b0;
      ways_3_metas_106_vld <= 1'b0;
      ways_3_metas_106_tag <= 51'h0;
      ways_3_metas_106_mru <= 1'b0;
      ways_3_metas_107_vld <= 1'b0;
      ways_3_metas_107_tag <= 51'h0;
      ways_3_metas_107_mru <= 1'b0;
      ways_3_metas_108_vld <= 1'b0;
      ways_3_metas_108_tag <= 51'h0;
      ways_3_metas_108_mru <= 1'b0;
      ways_3_metas_109_vld <= 1'b0;
      ways_3_metas_109_tag <= 51'h0;
      ways_3_metas_109_mru <= 1'b0;
      ways_3_metas_110_vld <= 1'b0;
      ways_3_metas_110_tag <= 51'h0;
      ways_3_metas_110_mru <= 1'b0;
      ways_3_metas_111_vld <= 1'b0;
      ways_3_metas_111_tag <= 51'h0;
      ways_3_metas_111_mru <= 1'b0;
      ways_3_metas_112_vld <= 1'b0;
      ways_3_metas_112_tag <= 51'h0;
      ways_3_metas_112_mru <= 1'b0;
      ways_3_metas_113_vld <= 1'b0;
      ways_3_metas_113_tag <= 51'h0;
      ways_3_metas_113_mru <= 1'b0;
      ways_3_metas_114_vld <= 1'b0;
      ways_3_metas_114_tag <= 51'h0;
      ways_3_metas_114_mru <= 1'b0;
      ways_3_metas_115_vld <= 1'b0;
      ways_3_metas_115_tag <= 51'h0;
      ways_3_metas_115_mru <= 1'b0;
      ways_3_metas_116_vld <= 1'b0;
      ways_3_metas_116_tag <= 51'h0;
      ways_3_metas_116_mru <= 1'b0;
      ways_3_metas_117_vld <= 1'b0;
      ways_3_metas_117_tag <= 51'h0;
      ways_3_metas_117_mru <= 1'b0;
      ways_3_metas_118_vld <= 1'b0;
      ways_3_metas_118_tag <= 51'h0;
      ways_3_metas_118_mru <= 1'b0;
      ways_3_metas_119_vld <= 1'b0;
      ways_3_metas_119_tag <= 51'h0;
      ways_3_metas_119_mru <= 1'b0;
      ways_3_metas_120_vld <= 1'b0;
      ways_3_metas_120_tag <= 51'h0;
      ways_3_metas_120_mru <= 1'b0;
      ways_3_metas_121_vld <= 1'b0;
      ways_3_metas_121_tag <= 51'h0;
      ways_3_metas_121_mru <= 1'b0;
      ways_3_metas_122_vld <= 1'b0;
      ways_3_metas_122_tag <= 51'h0;
      ways_3_metas_122_mru <= 1'b0;
      ways_3_metas_123_vld <= 1'b0;
      ways_3_metas_123_tag <= 51'h0;
      ways_3_metas_123_mru <= 1'b0;
      ways_3_metas_124_vld <= 1'b0;
      ways_3_metas_124_tag <= 51'h0;
      ways_3_metas_124_mru <= 1'b0;
      ways_3_metas_125_vld <= 1'b0;
      ways_3_metas_125_tag <= 51'h0;
      ways_3_metas_125_mru <= 1'b0;
      ways_3_metas_126_vld <= 1'b0;
      ways_3_metas_126_tag <= 51'h0;
      ways_3_metas_126_mru <= 1'b0;
      ways_3_metas_127_vld <= 1'b0;
      ways_3_metas_127_tag <= 51'h0;
      ways_3_metas_127_mru <= 1'b0;
      flush_busy <= 1'b0;
      flush_cnt_value <= 7'h0;
      cpu_cmd_ready_1 <= 1'b1;
      next_level_cmd_valid_1 <= 1'b0;
      next_level_data_cnt_value <= 3'b000;
    end else begin
      flush_cnt_value <= flush_cnt_valueNext;
      next_level_data_cnt_value <= next_level_data_cnt_valueNext;
      if(when_DCache_l123) begin
        next_level_cmd_valid_1 <= 1'b1;
      end else begin
        next_level_cmd_valid_1 <= 1'b0;
      end
      if(flush) begin
        flush_busy <= 1'b1;
      end else begin
        if(flush_done) begin
          flush_busy <= 1'b0;
        end
      end
      if(flush_busy) begin
        if(_zz_131) begin
          ways_0_metas_0_mru <= 1'b0;
        end
        if(_zz_132) begin
          ways_0_metas_1_mru <= 1'b0;
        end
        if(_zz_133) begin
          ways_0_metas_2_mru <= 1'b0;
        end
        if(_zz_134) begin
          ways_0_metas_3_mru <= 1'b0;
        end
        if(_zz_135) begin
          ways_0_metas_4_mru <= 1'b0;
        end
        if(_zz_136) begin
          ways_0_metas_5_mru <= 1'b0;
        end
        if(_zz_137) begin
          ways_0_metas_6_mru <= 1'b0;
        end
        if(_zz_138) begin
          ways_0_metas_7_mru <= 1'b0;
        end
        if(_zz_139) begin
          ways_0_metas_8_mru <= 1'b0;
        end
        if(_zz_140) begin
          ways_0_metas_9_mru <= 1'b0;
        end
        if(_zz_141) begin
          ways_0_metas_10_mru <= 1'b0;
        end
        if(_zz_142) begin
          ways_0_metas_11_mru <= 1'b0;
        end
        if(_zz_143) begin
          ways_0_metas_12_mru <= 1'b0;
        end
        if(_zz_144) begin
          ways_0_metas_13_mru <= 1'b0;
        end
        if(_zz_145) begin
          ways_0_metas_14_mru <= 1'b0;
        end
        if(_zz_146) begin
          ways_0_metas_15_mru <= 1'b0;
        end
        if(_zz_147) begin
          ways_0_metas_16_mru <= 1'b0;
        end
        if(_zz_148) begin
          ways_0_metas_17_mru <= 1'b0;
        end
        if(_zz_149) begin
          ways_0_metas_18_mru <= 1'b0;
        end
        if(_zz_150) begin
          ways_0_metas_19_mru <= 1'b0;
        end
        if(_zz_151) begin
          ways_0_metas_20_mru <= 1'b0;
        end
        if(_zz_152) begin
          ways_0_metas_21_mru <= 1'b0;
        end
        if(_zz_153) begin
          ways_0_metas_22_mru <= 1'b0;
        end
        if(_zz_154) begin
          ways_0_metas_23_mru <= 1'b0;
        end
        if(_zz_155) begin
          ways_0_metas_24_mru <= 1'b0;
        end
        if(_zz_156) begin
          ways_0_metas_25_mru <= 1'b0;
        end
        if(_zz_157) begin
          ways_0_metas_26_mru <= 1'b0;
        end
        if(_zz_158) begin
          ways_0_metas_27_mru <= 1'b0;
        end
        if(_zz_159) begin
          ways_0_metas_28_mru <= 1'b0;
        end
        if(_zz_160) begin
          ways_0_metas_29_mru <= 1'b0;
        end
        if(_zz_161) begin
          ways_0_metas_30_mru <= 1'b0;
        end
        if(_zz_162) begin
          ways_0_metas_31_mru <= 1'b0;
        end
        if(_zz_163) begin
          ways_0_metas_32_mru <= 1'b0;
        end
        if(_zz_164) begin
          ways_0_metas_33_mru <= 1'b0;
        end
        if(_zz_165) begin
          ways_0_metas_34_mru <= 1'b0;
        end
        if(_zz_166) begin
          ways_0_metas_35_mru <= 1'b0;
        end
        if(_zz_167) begin
          ways_0_metas_36_mru <= 1'b0;
        end
        if(_zz_168) begin
          ways_0_metas_37_mru <= 1'b0;
        end
        if(_zz_169) begin
          ways_0_metas_38_mru <= 1'b0;
        end
        if(_zz_170) begin
          ways_0_metas_39_mru <= 1'b0;
        end
        if(_zz_171) begin
          ways_0_metas_40_mru <= 1'b0;
        end
        if(_zz_172) begin
          ways_0_metas_41_mru <= 1'b0;
        end
        if(_zz_173) begin
          ways_0_metas_42_mru <= 1'b0;
        end
        if(_zz_174) begin
          ways_0_metas_43_mru <= 1'b0;
        end
        if(_zz_175) begin
          ways_0_metas_44_mru <= 1'b0;
        end
        if(_zz_176) begin
          ways_0_metas_45_mru <= 1'b0;
        end
        if(_zz_177) begin
          ways_0_metas_46_mru <= 1'b0;
        end
        if(_zz_178) begin
          ways_0_metas_47_mru <= 1'b0;
        end
        if(_zz_179) begin
          ways_0_metas_48_mru <= 1'b0;
        end
        if(_zz_180) begin
          ways_0_metas_49_mru <= 1'b0;
        end
        if(_zz_181) begin
          ways_0_metas_50_mru <= 1'b0;
        end
        if(_zz_182) begin
          ways_0_metas_51_mru <= 1'b0;
        end
        if(_zz_183) begin
          ways_0_metas_52_mru <= 1'b0;
        end
        if(_zz_184) begin
          ways_0_metas_53_mru <= 1'b0;
        end
        if(_zz_185) begin
          ways_0_metas_54_mru <= 1'b0;
        end
        if(_zz_186) begin
          ways_0_metas_55_mru <= 1'b0;
        end
        if(_zz_187) begin
          ways_0_metas_56_mru <= 1'b0;
        end
        if(_zz_188) begin
          ways_0_metas_57_mru <= 1'b0;
        end
        if(_zz_189) begin
          ways_0_metas_58_mru <= 1'b0;
        end
        if(_zz_190) begin
          ways_0_metas_59_mru <= 1'b0;
        end
        if(_zz_191) begin
          ways_0_metas_60_mru <= 1'b0;
        end
        if(_zz_192) begin
          ways_0_metas_61_mru <= 1'b0;
        end
        if(_zz_193) begin
          ways_0_metas_62_mru <= 1'b0;
        end
        if(_zz_194) begin
          ways_0_metas_63_mru <= 1'b0;
        end
        if(_zz_195) begin
          ways_0_metas_64_mru <= 1'b0;
        end
        if(_zz_196) begin
          ways_0_metas_65_mru <= 1'b0;
        end
        if(_zz_197) begin
          ways_0_metas_66_mru <= 1'b0;
        end
        if(_zz_198) begin
          ways_0_metas_67_mru <= 1'b0;
        end
        if(_zz_199) begin
          ways_0_metas_68_mru <= 1'b0;
        end
        if(_zz_200) begin
          ways_0_metas_69_mru <= 1'b0;
        end
        if(_zz_201) begin
          ways_0_metas_70_mru <= 1'b0;
        end
        if(_zz_202) begin
          ways_0_metas_71_mru <= 1'b0;
        end
        if(_zz_203) begin
          ways_0_metas_72_mru <= 1'b0;
        end
        if(_zz_204) begin
          ways_0_metas_73_mru <= 1'b0;
        end
        if(_zz_205) begin
          ways_0_metas_74_mru <= 1'b0;
        end
        if(_zz_206) begin
          ways_0_metas_75_mru <= 1'b0;
        end
        if(_zz_207) begin
          ways_0_metas_76_mru <= 1'b0;
        end
        if(_zz_208) begin
          ways_0_metas_77_mru <= 1'b0;
        end
        if(_zz_209) begin
          ways_0_metas_78_mru <= 1'b0;
        end
        if(_zz_210) begin
          ways_0_metas_79_mru <= 1'b0;
        end
        if(_zz_211) begin
          ways_0_metas_80_mru <= 1'b0;
        end
        if(_zz_212) begin
          ways_0_metas_81_mru <= 1'b0;
        end
        if(_zz_213) begin
          ways_0_metas_82_mru <= 1'b0;
        end
        if(_zz_214) begin
          ways_0_metas_83_mru <= 1'b0;
        end
        if(_zz_215) begin
          ways_0_metas_84_mru <= 1'b0;
        end
        if(_zz_216) begin
          ways_0_metas_85_mru <= 1'b0;
        end
        if(_zz_217) begin
          ways_0_metas_86_mru <= 1'b0;
        end
        if(_zz_218) begin
          ways_0_metas_87_mru <= 1'b0;
        end
        if(_zz_219) begin
          ways_0_metas_88_mru <= 1'b0;
        end
        if(_zz_220) begin
          ways_0_metas_89_mru <= 1'b0;
        end
        if(_zz_221) begin
          ways_0_metas_90_mru <= 1'b0;
        end
        if(_zz_222) begin
          ways_0_metas_91_mru <= 1'b0;
        end
        if(_zz_223) begin
          ways_0_metas_92_mru <= 1'b0;
        end
        if(_zz_224) begin
          ways_0_metas_93_mru <= 1'b0;
        end
        if(_zz_225) begin
          ways_0_metas_94_mru <= 1'b0;
        end
        if(_zz_226) begin
          ways_0_metas_95_mru <= 1'b0;
        end
        if(_zz_227) begin
          ways_0_metas_96_mru <= 1'b0;
        end
        if(_zz_228) begin
          ways_0_metas_97_mru <= 1'b0;
        end
        if(_zz_229) begin
          ways_0_metas_98_mru <= 1'b0;
        end
        if(_zz_230) begin
          ways_0_metas_99_mru <= 1'b0;
        end
        if(_zz_231) begin
          ways_0_metas_100_mru <= 1'b0;
        end
        if(_zz_232) begin
          ways_0_metas_101_mru <= 1'b0;
        end
        if(_zz_233) begin
          ways_0_metas_102_mru <= 1'b0;
        end
        if(_zz_234) begin
          ways_0_metas_103_mru <= 1'b0;
        end
        if(_zz_235) begin
          ways_0_metas_104_mru <= 1'b0;
        end
        if(_zz_236) begin
          ways_0_metas_105_mru <= 1'b0;
        end
        if(_zz_237) begin
          ways_0_metas_106_mru <= 1'b0;
        end
        if(_zz_238) begin
          ways_0_metas_107_mru <= 1'b0;
        end
        if(_zz_239) begin
          ways_0_metas_108_mru <= 1'b0;
        end
        if(_zz_240) begin
          ways_0_metas_109_mru <= 1'b0;
        end
        if(_zz_241) begin
          ways_0_metas_110_mru <= 1'b0;
        end
        if(_zz_242) begin
          ways_0_metas_111_mru <= 1'b0;
        end
        if(_zz_243) begin
          ways_0_metas_112_mru <= 1'b0;
        end
        if(_zz_244) begin
          ways_0_metas_113_mru <= 1'b0;
        end
        if(_zz_245) begin
          ways_0_metas_114_mru <= 1'b0;
        end
        if(_zz_246) begin
          ways_0_metas_115_mru <= 1'b0;
        end
        if(_zz_247) begin
          ways_0_metas_116_mru <= 1'b0;
        end
        if(_zz_248) begin
          ways_0_metas_117_mru <= 1'b0;
        end
        if(_zz_249) begin
          ways_0_metas_118_mru <= 1'b0;
        end
        if(_zz_250) begin
          ways_0_metas_119_mru <= 1'b0;
        end
        if(_zz_251) begin
          ways_0_metas_120_mru <= 1'b0;
        end
        if(_zz_252) begin
          ways_0_metas_121_mru <= 1'b0;
        end
        if(_zz_253) begin
          ways_0_metas_122_mru <= 1'b0;
        end
        if(_zz_254) begin
          ways_0_metas_123_mru <= 1'b0;
        end
        if(_zz_255) begin
          ways_0_metas_124_mru <= 1'b0;
        end
        if(_zz_256) begin
          ways_0_metas_125_mru <= 1'b0;
        end
        if(_zz_257) begin
          ways_0_metas_126_mru <= 1'b0;
        end
        if(_zz_258) begin
          ways_0_metas_127_mru <= 1'b0;
        end
        if(_zz_131) begin
          ways_0_metas_0_vld <= 1'b0;
        end
        if(_zz_132) begin
          ways_0_metas_1_vld <= 1'b0;
        end
        if(_zz_133) begin
          ways_0_metas_2_vld <= 1'b0;
        end
        if(_zz_134) begin
          ways_0_metas_3_vld <= 1'b0;
        end
        if(_zz_135) begin
          ways_0_metas_4_vld <= 1'b0;
        end
        if(_zz_136) begin
          ways_0_metas_5_vld <= 1'b0;
        end
        if(_zz_137) begin
          ways_0_metas_6_vld <= 1'b0;
        end
        if(_zz_138) begin
          ways_0_metas_7_vld <= 1'b0;
        end
        if(_zz_139) begin
          ways_0_metas_8_vld <= 1'b0;
        end
        if(_zz_140) begin
          ways_0_metas_9_vld <= 1'b0;
        end
        if(_zz_141) begin
          ways_0_metas_10_vld <= 1'b0;
        end
        if(_zz_142) begin
          ways_0_metas_11_vld <= 1'b0;
        end
        if(_zz_143) begin
          ways_0_metas_12_vld <= 1'b0;
        end
        if(_zz_144) begin
          ways_0_metas_13_vld <= 1'b0;
        end
        if(_zz_145) begin
          ways_0_metas_14_vld <= 1'b0;
        end
        if(_zz_146) begin
          ways_0_metas_15_vld <= 1'b0;
        end
        if(_zz_147) begin
          ways_0_metas_16_vld <= 1'b0;
        end
        if(_zz_148) begin
          ways_0_metas_17_vld <= 1'b0;
        end
        if(_zz_149) begin
          ways_0_metas_18_vld <= 1'b0;
        end
        if(_zz_150) begin
          ways_0_metas_19_vld <= 1'b0;
        end
        if(_zz_151) begin
          ways_0_metas_20_vld <= 1'b0;
        end
        if(_zz_152) begin
          ways_0_metas_21_vld <= 1'b0;
        end
        if(_zz_153) begin
          ways_0_metas_22_vld <= 1'b0;
        end
        if(_zz_154) begin
          ways_0_metas_23_vld <= 1'b0;
        end
        if(_zz_155) begin
          ways_0_metas_24_vld <= 1'b0;
        end
        if(_zz_156) begin
          ways_0_metas_25_vld <= 1'b0;
        end
        if(_zz_157) begin
          ways_0_metas_26_vld <= 1'b0;
        end
        if(_zz_158) begin
          ways_0_metas_27_vld <= 1'b0;
        end
        if(_zz_159) begin
          ways_0_metas_28_vld <= 1'b0;
        end
        if(_zz_160) begin
          ways_0_metas_29_vld <= 1'b0;
        end
        if(_zz_161) begin
          ways_0_metas_30_vld <= 1'b0;
        end
        if(_zz_162) begin
          ways_0_metas_31_vld <= 1'b0;
        end
        if(_zz_163) begin
          ways_0_metas_32_vld <= 1'b0;
        end
        if(_zz_164) begin
          ways_0_metas_33_vld <= 1'b0;
        end
        if(_zz_165) begin
          ways_0_metas_34_vld <= 1'b0;
        end
        if(_zz_166) begin
          ways_0_metas_35_vld <= 1'b0;
        end
        if(_zz_167) begin
          ways_0_metas_36_vld <= 1'b0;
        end
        if(_zz_168) begin
          ways_0_metas_37_vld <= 1'b0;
        end
        if(_zz_169) begin
          ways_0_metas_38_vld <= 1'b0;
        end
        if(_zz_170) begin
          ways_0_metas_39_vld <= 1'b0;
        end
        if(_zz_171) begin
          ways_0_metas_40_vld <= 1'b0;
        end
        if(_zz_172) begin
          ways_0_metas_41_vld <= 1'b0;
        end
        if(_zz_173) begin
          ways_0_metas_42_vld <= 1'b0;
        end
        if(_zz_174) begin
          ways_0_metas_43_vld <= 1'b0;
        end
        if(_zz_175) begin
          ways_0_metas_44_vld <= 1'b0;
        end
        if(_zz_176) begin
          ways_0_metas_45_vld <= 1'b0;
        end
        if(_zz_177) begin
          ways_0_metas_46_vld <= 1'b0;
        end
        if(_zz_178) begin
          ways_0_metas_47_vld <= 1'b0;
        end
        if(_zz_179) begin
          ways_0_metas_48_vld <= 1'b0;
        end
        if(_zz_180) begin
          ways_0_metas_49_vld <= 1'b0;
        end
        if(_zz_181) begin
          ways_0_metas_50_vld <= 1'b0;
        end
        if(_zz_182) begin
          ways_0_metas_51_vld <= 1'b0;
        end
        if(_zz_183) begin
          ways_0_metas_52_vld <= 1'b0;
        end
        if(_zz_184) begin
          ways_0_metas_53_vld <= 1'b0;
        end
        if(_zz_185) begin
          ways_0_metas_54_vld <= 1'b0;
        end
        if(_zz_186) begin
          ways_0_metas_55_vld <= 1'b0;
        end
        if(_zz_187) begin
          ways_0_metas_56_vld <= 1'b0;
        end
        if(_zz_188) begin
          ways_0_metas_57_vld <= 1'b0;
        end
        if(_zz_189) begin
          ways_0_metas_58_vld <= 1'b0;
        end
        if(_zz_190) begin
          ways_0_metas_59_vld <= 1'b0;
        end
        if(_zz_191) begin
          ways_0_metas_60_vld <= 1'b0;
        end
        if(_zz_192) begin
          ways_0_metas_61_vld <= 1'b0;
        end
        if(_zz_193) begin
          ways_0_metas_62_vld <= 1'b0;
        end
        if(_zz_194) begin
          ways_0_metas_63_vld <= 1'b0;
        end
        if(_zz_195) begin
          ways_0_metas_64_vld <= 1'b0;
        end
        if(_zz_196) begin
          ways_0_metas_65_vld <= 1'b0;
        end
        if(_zz_197) begin
          ways_0_metas_66_vld <= 1'b0;
        end
        if(_zz_198) begin
          ways_0_metas_67_vld <= 1'b0;
        end
        if(_zz_199) begin
          ways_0_metas_68_vld <= 1'b0;
        end
        if(_zz_200) begin
          ways_0_metas_69_vld <= 1'b0;
        end
        if(_zz_201) begin
          ways_0_metas_70_vld <= 1'b0;
        end
        if(_zz_202) begin
          ways_0_metas_71_vld <= 1'b0;
        end
        if(_zz_203) begin
          ways_0_metas_72_vld <= 1'b0;
        end
        if(_zz_204) begin
          ways_0_metas_73_vld <= 1'b0;
        end
        if(_zz_205) begin
          ways_0_metas_74_vld <= 1'b0;
        end
        if(_zz_206) begin
          ways_0_metas_75_vld <= 1'b0;
        end
        if(_zz_207) begin
          ways_0_metas_76_vld <= 1'b0;
        end
        if(_zz_208) begin
          ways_0_metas_77_vld <= 1'b0;
        end
        if(_zz_209) begin
          ways_0_metas_78_vld <= 1'b0;
        end
        if(_zz_210) begin
          ways_0_metas_79_vld <= 1'b0;
        end
        if(_zz_211) begin
          ways_0_metas_80_vld <= 1'b0;
        end
        if(_zz_212) begin
          ways_0_metas_81_vld <= 1'b0;
        end
        if(_zz_213) begin
          ways_0_metas_82_vld <= 1'b0;
        end
        if(_zz_214) begin
          ways_0_metas_83_vld <= 1'b0;
        end
        if(_zz_215) begin
          ways_0_metas_84_vld <= 1'b0;
        end
        if(_zz_216) begin
          ways_0_metas_85_vld <= 1'b0;
        end
        if(_zz_217) begin
          ways_0_metas_86_vld <= 1'b0;
        end
        if(_zz_218) begin
          ways_0_metas_87_vld <= 1'b0;
        end
        if(_zz_219) begin
          ways_0_metas_88_vld <= 1'b0;
        end
        if(_zz_220) begin
          ways_0_metas_89_vld <= 1'b0;
        end
        if(_zz_221) begin
          ways_0_metas_90_vld <= 1'b0;
        end
        if(_zz_222) begin
          ways_0_metas_91_vld <= 1'b0;
        end
        if(_zz_223) begin
          ways_0_metas_92_vld <= 1'b0;
        end
        if(_zz_224) begin
          ways_0_metas_93_vld <= 1'b0;
        end
        if(_zz_225) begin
          ways_0_metas_94_vld <= 1'b0;
        end
        if(_zz_226) begin
          ways_0_metas_95_vld <= 1'b0;
        end
        if(_zz_227) begin
          ways_0_metas_96_vld <= 1'b0;
        end
        if(_zz_228) begin
          ways_0_metas_97_vld <= 1'b0;
        end
        if(_zz_229) begin
          ways_0_metas_98_vld <= 1'b0;
        end
        if(_zz_230) begin
          ways_0_metas_99_vld <= 1'b0;
        end
        if(_zz_231) begin
          ways_0_metas_100_vld <= 1'b0;
        end
        if(_zz_232) begin
          ways_0_metas_101_vld <= 1'b0;
        end
        if(_zz_233) begin
          ways_0_metas_102_vld <= 1'b0;
        end
        if(_zz_234) begin
          ways_0_metas_103_vld <= 1'b0;
        end
        if(_zz_235) begin
          ways_0_metas_104_vld <= 1'b0;
        end
        if(_zz_236) begin
          ways_0_metas_105_vld <= 1'b0;
        end
        if(_zz_237) begin
          ways_0_metas_106_vld <= 1'b0;
        end
        if(_zz_238) begin
          ways_0_metas_107_vld <= 1'b0;
        end
        if(_zz_239) begin
          ways_0_metas_108_vld <= 1'b0;
        end
        if(_zz_240) begin
          ways_0_metas_109_vld <= 1'b0;
        end
        if(_zz_241) begin
          ways_0_metas_110_vld <= 1'b0;
        end
        if(_zz_242) begin
          ways_0_metas_111_vld <= 1'b0;
        end
        if(_zz_243) begin
          ways_0_metas_112_vld <= 1'b0;
        end
        if(_zz_244) begin
          ways_0_metas_113_vld <= 1'b0;
        end
        if(_zz_245) begin
          ways_0_metas_114_vld <= 1'b0;
        end
        if(_zz_246) begin
          ways_0_metas_115_vld <= 1'b0;
        end
        if(_zz_247) begin
          ways_0_metas_116_vld <= 1'b0;
        end
        if(_zz_248) begin
          ways_0_metas_117_vld <= 1'b0;
        end
        if(_zz_249) begin
          ways_0_metas_118_vld <= 1'b0;
        end
        if(_zz_250) begin
          ways_0_metas_119_vld <= 1'b0;
        end
        if(_zz_251) begin
          ways_0_metas_120_vld <= 1'b0;
        end
        if(_zz_252) begin
          ways_0_metas_121_vld <= 1'b0;
        end
        if(_zz_253) begin
          ways_0_metas_122_vld <= 1'b0;
        end
        if(_zz_254) begin
          ways_0_metas_123_vld <= 1'b0;
        end
        if(_zz_255) begin
          ways_0_metas_124_vld <= 1'b0;
        end
        if(_zz_256) begin
          ways_0_metas_125_vld <= 1'b0;
        end
        if(_zz_257) begin
          ways_0_metas_126_vld <= 1'b0;
        end
        if(_zz_258) begin
          ways_0_metas_127_vld <= 1'b0;
        end
      end else begin
        if(when_DCache_l217) begin
          if(cache_hit_0) begin
            if(_zz_2) begin
              ways_0_metas_0_mru <= 1'b1;
            end
            if(_zz_3) begin
              ways_0_metas_1_mru <= 1'b1;
            end
            if(_zz_4) begin
              ways_0_metas_2_mru <= 1'b1;
            end
            if(_zz_5) begin
              ways_0_metas_3_mru <= 1'b1;
            end
            if(_zz_6) begin
              ways_0_metas_4_mru <= 1'b1;
            end
            if(_zz_7) begin
              ways_0_metas_5_mru <= 1'b1;
            end
            if(_zz_8) begin
              ways_0_metas_6_mru <= 1'b1;
            end
            if(_zz_9) begin
              ways_0_metas_7_mru <= 1'b1;
            end
            if(_zz_10) begin
              ways_0_metas_8_mru <= 1'b1;
            end
            if(_zz_11) begin
              ways_0_metas_9_mru <= 1'b1;
            end
            if(_zz_12) begin
              ways_0_metas_10_mru <= 1'b1;
            end
            if(_zz_13) begin
              ways_0_metas_11_mru <= 1'b1;
            end
            if(_zz_14) begin
              ways_0_metas_12_mru <= 1'b1;
            end
            if(_zz_15) begin
              ways_0_metas_13_mru <= 1'b1;
            end
            if(_zz_16) begin
              ways_0_metas_14_mru <= 1'b1;
            end
            if(_zz_17) begin
              ways_0_metas_15_mru <= 1'b1;
            end
            if(_zz_18) begin
              ways_0_metas_16_mru <= 1'b1;
            end
            if(_zz_19) begin
              ways_0_metas_17_mru <= 1'b1;
            end
            if(_zz_20) begin
              ways_0_metas_18_mru <= 1'b1;
            end
            if(_zz_21) begin
              ways_0_metas_19_mru <= 1'b1;
            end
            if(_zz_22) begin
              ways_0_metas_20_mru <= 1'b1;
            end
            if(_zz_23) begin
              ways_0_metas_21_mru <= 1'b1;
            end
            if(_zz_24) begin
              ways_0_metas_22_mru <= 1'b1;
            end
            if(_zz_25) begin
              ways_0_metas_23_mru <= 1'b1;
            end
            if(_zz_26) begin
              ways_0_metas_24_mru <= 1'b1;
            end
            if(_zz_27) begin
              ways_0_metas_25_mru <= 1'b1;
            end
            if(_zz_28) begin
              ways_0_metas_26_mru <= 1'b1;
            end
            if(_zz_29) begin
              ways_0_metas_27_mru <= 1'b1;
            end
            if(_zz_30) begin
              ways_0_metas_28_mru <= 1'b1;
            end
            if(_zz_31) begin
              ways_0_metas_29_mru <= 1'b1;
            end
            if(_zz_32) begin
              ways_0_metas_30_mru <= 1'b1;
            end
            if(_zz_33) begin
              ways_0_metas_31_mru <= 1'b1;
            end
            if(_zz_34) begin
              ways_0_metas_32_mru <= 1'b1;
            end
            if(_zz_35) begin
              ways_0_metas_33_mru <= 1'b1;
            end
            if(_zz_36) begin
              ways_0_metas_34_mru <= 1'b1;
            end
            if(_zz_37) begin
              ways_0_metas_35_mru <= 1'b1;
            end
            if(_zz_38) begin
              ways_0_metas_36_mru <= 1'b1;
            end
            if(_zz_39) begin
              ways_0_metas_37_mru <= 1'b1;
            end
            if(_zz_40) begin
              ways_0_metas_38_mru <= 1'b1;
            end
            if(_zz_41) begin
              ways_0_metas_39_mru <= 1'b1;
            end
            if(_zz_42) begin
              ways_0_metas_40_mru <= 1'b1;
            end
            if(_zz_43) begin
              ways_0_metas_41_mru <= 1'b1;
            end
            if(_zz_44) begin
              ways_0_metas_42_mru <= 1'b1;
            end
            if(_zz_45) begin
              ways_0_metas_43_mru <= 1'b1;
            end
            if(_zz_46) begin
              ways_0_metas_44_mru <= 1'b1;
            end
            if(_zz_47) begin
              ways_0_metas_45_mru <= 1'b1;
            end
            if(_zz_48) begin
              ways_0_metas_46_mru <= 1'b1;
            end
            if(_zz_49) begin
              ways_0_metas_47_mru <= 1'b1;
            end
            if(_zz_50) begin
              ways_0_metas_48_mru <= 1'b1;
            end
            if(_zz_51) begin
              ways_0_metas_49_mru <= 1'b1;
            end
            if(_zz_52) begin
              ways_0_metas_50_mru <= 1'b1;
            end
            if(_zz_53) begin
              ways_0_metas_51_mru <= 1'b1;
            end
            if(_zz_54) begin
              ways_0_metas_52_mru <= 1'b1;
            end
            if(_zz_55) begin
              ways_0_metas_53_mru <= 1'b1;
            end
            if(_zz_56) begin
              ways_0_metas_54_mru <= 1'b1;
            end
            if(_zz_57) begin
              ways_0_metas_55_mru <= 1'b1;
            end
            if(_zz_58) begin
              ways_0_metas_56_mru <= 1'b1;
            end
            if(_zz_59) begin
              ways_0_metas_57_mru <= 1'b1;
            end
            if(_zz_60) begin
              ways_0_metas_58_mru <= 1'b1;
            end
            if(_zz_61) begin
              ways_0_metas_59_mru <= 1'b1;
            end
            if(_zz_62) begin
              ways_0_metas_60_mru <= 1'b1;
            end
            if(_zz_63) begin
              ways_0_metas_61_mru <= 1'b1;
            end
            if(_zz_64) begin
              ways_0_metas_62_mru <= 1'b1;
            end
            if(_zz_65) begin
              ways_0_metas_63_mru <= 1'b1;
            end
            if(_zz_66) begin
              ways_0_metas_64_mru <= 1'b1;
            end
            if(_zz_67) begin
              ways_0_metas_65_mru <= 1'b1;
            end
            if(_zz_68) begin
              ways_0_metas_66_mru <= 1'b1;
            end
            if(_zz_69) begin
              ways_0_metas_67_mru <= 1'b1;
            end
            if(_zz_70) begin
              ways_0_metas_68_mru <= 1'b1;
            end
            if(_zz_71) begin
              ways_0_metas_69_mru <= 1'b1;
            end
            if(_zz_72) begin
              ways_0_metas_70_mru <= 1'b1;
            end
            if(_zz_73) begin
              ways_0_metas_71_mru <= 1'b1;
            end
            if(_zz_74) begin
              ways_0_metas_72_mru <= 1'b1;
            end
            if(_zz_75) begin
              ways_0_metas_73_mru <= 1'b1;
            end
            if(_zz_76) begin
              ways_0_metas_74_mru <= 1'b1;
            end
            if(_zz_77) begin
              ways_0_metas_75_mru <= 1'b1;
            end
            if(_zz_78) begin
              ways_0_metas_76_mru <= 1'b1;
            end
            if(_zz_79) begin
              ways_0_metas_77_mru <= 1'b1;
            end
            if(_zz_80) begin
              ways_0_metas_78_mru <= 1'b1;
            end
            if(_zz_81) begin
              ways_0_metas_79_mru <= 1'b1;
            end
            if(_zz_82) begin
              ways_0_metas_80_mru <= 1'b1;
            end
            if(_zz_83) begin
              ways_0_metas_81_mru <= 1'b1;
            end
            if(_zz_84) begin
              ways_0_metas_82_mru <= 1'b1;
            end
            if(_zz_85) begin
              ways_0_metas_83_mru <= 1'b1;
            end
            if(_zz_86) begin
              ways_0_metas_84_mru <= 1'b1;
            end
            if(_zz_87) begin
              ways_0_metas_85_mru <= 1'b1;
            end
            if(_zz_88) begin
              ways_0_metas_86_mru <= 1'b1;
            end
            if(_zz_89) begin
              ways_0_metas_87_mru <= 1'b1;
            end
            if(_zz_90) begin
              ways_0_metas_88_mru <= 1'b1;
            end
            if(_zz_91) begin
              ways_0_metas_89_mru <= 1'b1;
            end
            if(_zz_92) begin
              ways_0_metas_90_mru <= 1'b1;
            end
            if(_zz_93) begin
              ways_0_metas_91_mru <= 1'b1;
            end
            if(_zz_94) begin
              ways_0_metas_92_mru <= 1'b1;
            end
            if(_zz_95) begin
              ways_0_metas_93_mru <= 1'b1;
            end
            if(_zz_96) begin
              ways_0_metas_94_mru <= 1'b1;
            end
            if(_zz_97) begin
              ways_0_metas_95_mru <= 1'b1;
            end
            if(_zz_98) begin
              ways_0_metas_96_mru <= 1'b1;
            end
            if(_zz_99) begin
              ways_0_metas_97_mru <= 1'b1;
            end
            if(_zz_100) begin
              ways_0_metas_98_mru <= 1'b1;
            end
            if(_zz_101) begin
              ways_0_metas_99_mru <= 1'b1;
            end
            if(_zz_102) begin
              ways_0_metas_100_mru <= 1'b1;
            end
            if(_zz_103) begin
              ways_0_metas_101_mru <= 1'b1;
            end
            if(_zz_104) begin
              ways_0_metas_102_mru <= 1'b1;
            end
            if(_zz_105) begin
              ways_0_metas_103_mru <= 1'b1;
            end
            if(_zz_106) begin
              ways_0_metas_104_mru <= 1'b1;
            end
            if(_zz_107) begin
              ways_0_metas_105_mru <= 1'b1;
            end
            if(_zz_108) begin
              ways_0_metas_106_mru <= 1'b1;
            end
            if(_zz_109) begin
              ways_0_metas_107_mru <= 1'b1;
            end
            if(_zz_110) begin
              ways_0_metas_108_mru <= 1'b1;
            end
            if(_zz_111) begin
              ways_0_metas_109_mru <= 1'b1;
            end
            if(_zz_112) begin
              ways_0_metas_110_mru <= 1'b1;
            end
            if(_zz_113) begin
              ways_0_metas_111_mru <= 1'b1;
            end
            if(_zz_114) begin
              ways_0_metas_112_mru <= 1'b1;
            end
            if(_zz_115) begin
              ways_0_metas_113_mru <= 1'b1;
            end
            if(_zz_116) begin
              ways_0_metas_114_mru <= 1'b1;
            end
            if(_zz_117) begin
              ways_0_metas_115_mru <= 1'b1;
            end
            if(_zz_118) begin
              ways_0_metas_116_mru <= 1'b1;
            end
            if(_zz_119) begin
              ways_0_metas_117_mru <= 1'b1;
            end
            if(_zz_120) begin
              ways_0_metas_118_mru <= 1'b1;
            end
            if(_zz_121) begin
              ways_0_metas_119_mru <= 1'b1;
            end
            if(_zz_122) begin
              ways_0_metas_120_mru <= 1'b1;
            end
            if(_zz_123) begin
              ways_0_metas_121_mru <= 1'b1;
            end
            if(_zz_124) begin
              ways_0_metas_122_mru <= 1'b1;
            end
            if(_zz_125) begin
              ways_0_metas_123_mru <= 1'b1;
            end
            if(_zz_126) begin
              ways_0_metas_124_mru <= 1'b1;
            end
            if(_zz_127) begin
              ways_0_metas_125_mru <= 1'b1;
            end
            if(_zz_128) begin
              ways_0_metas_126_mru <= 1'b1;
            end
            if(_zz_129) begin
              ways_0_metas_127_mru <= 1'b1;
            end
          end else begin
            if(_zz_2) begin
              ways_0_metas_0_mru <= 1'b0;
            end
            if(_zz_3) begin
              ways_0_metas_1_mru <= 1'b0;
            end
            if(_zz_4) begin
              ways_0_metas_2_mru <= 1'b0;
            end
            if(_zz_5) begin
              ways_0_metas_3_mru <= 1'b0;
            end
            if(_zz_6) begin
              ways_0_metas_4_mru <= 1'b0;
            end
            if(_zz_7) begin
              ways_0_metas_5_mru <= 1'b0;
            end
            if(_zz_8) begin
              ways_0_metas_6_mru <= 1'b0;
            end
            if(_zz_9) begin
              ways_0_metas_7_mru <= 1'b0;
            end
            if(_zz_10) begin
              ways_0_metas_8_mru <= 1'b0;
            end
            if(_zz_11) begin
              ways_0_metas_9_mru <= 1'b0;
            end
            if(_zz_12) begin
              ways_0_metas_10_mru <= 1'b0;
            end
            if(_zz_13) begin
              ways_0_metas_11_mru <= 1'b0;
            end
            if(_zz_14) begin
              ways_0_metas_12_mru <= 1'b0;
            end
            if(_zz_15) begin
              ways_0_metas_13_mru <= 1'b0;
            end
            if(_zz_16) begin
              ways_0_metas_14_mru <= 1'b0;
            end
            if(_zz_17) begin
              ways_0_metas_15_mru <= 1'b0;
            end
            if(_zz_18) begin
              ways_0_metas_16_mru <= 1'b0;
            end
            if(_zz_19) begin
              ways_0_metas_17_mru <= 1'b0;
            end
            if(_zz_20) begin
              ways_0_metas_18_mru <= 1'b0;
            end
            if(_zz_21) begin
              ways_0_metas_19_mru <= 1'b0;
            end
            if(_zz_22) begin
              ways_0_metas_20_mru <= 1'b0;
            end
            if(_zz_23) begin
              ways_0_metas_21_mru <= 1'b0;
            end
            if(_zz_24) begin
              ways_0_metas_22_mru <= 1'b0;
            end
            if(_zz_25) begin
              ways_0_metas_23_mru <= 1'b0;
            end
            if(_zz_26) begin
              ways_0_metas_24_mru <= 1'b0;
            end
            if(_zz_27) begin
              ways_0_metas_25_mru <= 1'b0;
            end
            if(_zz_28) begin
              ways_0_metas_26_mru <= 1'b0;
            end
            if(_zz_29) begin
              ways_0_metas_27_mru <= 1'b0;
            end
            if(_zz_30) begin
              ways_0_metas_28_mru <= 1'b0;
            end
            if(_zz_31) begin
              ways_0_metas_29_mru <= 1'b0;
            end
            if(_zz_32) begin
              ways_0_metas_30_mru <= 1'b0;
            end
            if(_zz_33) begin
              ways_0_metas_31_mru <= 1'b0;
            end
            if(_zz_34) begin
              ways_0_metas_32_mru <= 1'b0;
            end
            if(_zz_35) begin
              ways_0_metas_33_mru <= 1'b0;
            end
            if(_zz_36) begin
              ways_0_metas_34_mru <= 1'b0;
            end
            if(_zz_37) begin
              ways_0_metas_35_mru <= 1'b0;
            end
            if(_zz_38) begin
              ways_0_metas_36_mru <= 1'b0;
            end
            if(_zz_39) begin
              ways_0_metas_37_mru <= 1'b0;
            end
            if(_zz_40) begin
              ways_0_metas_38_mru <= 1'b0;
            end
            if(_zz_41) begin
              ways_0_metas_39_mru <= 1'b0;
            end
            if(_zz_42) begin
              ways_0_metas_40_mru <= 1'b0;
            end
            if(_zz_43) begin
              ways_0_metas_41_mru <= 1'b0;
            end
            if(_zz_44) begin
              ways_0_metas_42_mru <= 1'b0;
            end
            if(_zz_45) begin
              ways_0_metas_43_mru <= 1'b0;
            end
            if(_zz_46) begin
              ways_0_metas_44_mru <= 1'b0;
            end
            if(_zz_47) begin
              ways_0_metas_45_mru <= 1'b0;
            end
            if(_zz_48) begin
              ways_0_metas_46_mru <= 1'b0;
            end
            if(_zz_49) begin
              ways_0_metas_47_mru <= 1'b0;
            end
            if(_zz_50) begin
              ways_0_metas_48_mru <= 1'b0;
            end
            if(_zz_51) begin
              ways_0_metas_49_mru <= 1'b0;
            end
            if(_zz_52) begin
              ways_0_metas_50_mru <= 1'b0;
            end
            if(_zz_53) begin
              ways_0_metas_51_mru <= 1'b0;
            end
            if(_zz_54) begin
              ways_0_metas_52_mru <= 1'b0;
            end
            if(_zz_55) begin
              ways_0_metas_53_mru <= 1'b0;
            end
            if(_zz_56) begin
              ways_0_metas_54_mru <= 1'b0;
            end
            if(_zz_57) begin
              ways_0_metas_55_mru <= 1'b0;
            end
            if(_zz_58) begin
              ways_0_metas_56_mru <= 1'b0;
            end
            if(_zz_59) begin
              ways_0_metas_57_mru <= 1'b0;
            end
            if(_zz_60) begin
              ways_0_metas_58_mru <= 1'b0;
            end
            if(_zz_61) begin
              ways_0_metas_59_mru <= 1'b0;
            end
            if(_zz_62) begin
              ways_0_metas_60_mru <= 1'b0;
            end
            if(_zz_63) begin
              ways_0_metas_61_mru <= 1'b0;
            end
            if(_zz_64) begin
              ways_0_metas_62_mru <= 1'b0;
            end
            if(_zz_65) begin
              ways_0_metas_63_mru <= 1'b0;
            end
            if(_zz_66) begin
              ways_0_metas_64_mru <= 1'b0;
            end
            if(_zz_67) begin
              ways_0_metas_65_mru <= 1'b0;
            end
            if(_zz_68) begin
              ways_0_metas_66_mru <= 1'b0;
            end
            if(_zz_69) begin
              ways_0_metas_67_mru <= 1'b0;
            end
            if(_zz_70) begin
              ways_0_metas_68_mru <= 1'b0;
            end
            if(_zz_71) begin
              ways_0_metas_69_mru <= 1'b0;
            end
            if(_zz_72) begin
              ways_0_metas_70_mru <= 1'b0;
            end
            if(_zz_73) begin
              ways_0_metas_71_mru <= 1'b0;
            end
            if(_zz_74) begin
              ways_0_metas_72_mru <= 1'b0;
            end
            if(_zz_75) begin
              ways_0_metas_73_mru <= 1'b0;
            end
            if(_zz_76) begin
              ways_0_metas_74_mru <= 1'b0;
            end
            if(_zz_77) begin
              ways_0_metas_75_mru <= 1'b0;
            end
            if(_zz_78) begin
              ways_0_metas_76_mru <= 1'b0;
            end
            if(_zz_79) begin
              ways_0_metas_77_mru <= 1'b0;
            end
            if(_zz_80) begin
              ways_0_metas_78_mru <= 1'b0;
            end
            if(_zz_81) begin
              ways_0_metas_79_mru <= 1'b0;
            end
            if(_zz_82) begin
              ways_0_metas_80_mru <= 1'b0;
            end
            if(_zz_83) begin
              ways_0_metas_81_mru <= 1'b0;
            end
            if(_zz_84) begin
              ways_0_metas_82_mru <= 1'b0;
            end
            if(_zz_85) begin
              ways_0_metas_83_mru <= 1'b0;
            end
            if(_zz_86) begin
              ways_0_metas_84_mru <= 1'b0;
            end
            if(_zz_87) begin
              ways_0_metas_85_mru <= 1'b0;
            end
            if(_zz_88) begin
              ways_0_metas_86_mru <= 1'b0;
            end
            if(_zz_89) begin
              ways_0_metas_87_mru <= 1'b0;
            end
            if(_zz_90) begin
              ways_0_metas_88_mru <= 1'b0;
            end
            if(_zz_91) begin
              ways_0_metas_89_mru <= 1'b0;
            end
            if(_zz_92) begin
              ways_0_metas_90_mru <= 1'b0;
            end
            if(_zz_93) begin
              ways_0_metas_91_mru <= 1'b0;
            end
            if(_zz_94) begin
              ways_0_metas_92_mru <= 1'b0;
            end
            if(_zz_95) begin
              ways_0_metas_93_mru <= 1'b0;
            end
            if(_zz_96) begin
              ways_0_metas_94_mru <= 1'b0;
            end
            if(_zz_97) begin
              ways_0_metas_95_mru <= 1'b0;
            end
            if(_zz_98) begin
              ways_0_metas_96_mru <= 1'b0;
            end
            if(_zz_99) begin
              ways_0_metas_97_mru <= 1'b0;
            end
            if(_zz_100) begin
              ways_0_metas_98_mru <= 1'b0;
            end
            if(_zz_101) begin
              ways_0_metas_99_mru <= 1'b0;
            end
            if(_zz_102) begin
              ways_0_metas_100_mru <= 1'b0;
            end
            if(_zz_103) begin
              ways_0_metas_101_mru <= 1'b0;
            end
            if(_zz_104) begin
              ways_0_metas_102_mru <= 1'b0;
            end
            if(_zz_105) begin
              ways_0_metas_103_mru <= 1'b0;
            end
            if(_zz_106) begin
              ways_0_metas_104_mru <= 1'b0;
            end
            if(_zz_107) begin
              ways_0_metas_105_mru <= 1'b0;
            end
            if(_zz_108) begin
              ways_0_metas_106_mru <= 1'b0;
            end
            if(_zz_109) begin
              ways_0_metas_107_mru <= 1'b0;
            end
            if(_zz_110) begin
              ways_0_metas_108_mru <= 1'b0;
            end
            if(_zz_111) begin
              ways_0_metas_109_mru <= 1'b0;
            end
            if(_zz_112) begin
              ways_0_metas_110_mru <= 1'b0;
            end
            if(_zz_113) begin
              ways_0_metas_111_mru <= 1'b0;
            end
            if(_zz_114) begin
              ways_0_metas_112_mru <= 1'b0;
            end
            if(_zz_115) begin
              ways_0_metas_113_mru <= 1'b0;
            end
            if(_zz_116) begin
              ways_0_metas_114_mru <= 1'b0;
            end
            if(_zz_117) begin
              ways_0_metas_115_mru <= 1'b0;
            end
            if(_zz_118) begin
              ways_0_metas_116_mru <= 1'b0;
            end
            if(_zz_119) begin
              ways_0_metas_117_mru <= 1'b0;
            end
            if(_zz_120) begin
              ways_0_metas_118_mru <= 1'b0;
            end
            if(_zz_121) begin
              ways_0_metas_119_mru <= 1'b0;
            end
            if(_zz_122) begin
              ways_0_metas_120_mru <= 1'b0;
            end
            if(_zz_123) begin
              ways_0_metas_121_mru <= 1'b0;
            end
            if(_zz_124) begin
              ways_0_metas_122_mru <= 1'b0;
            end
            if(_zz_125) begin
              ways_0_metas_123_mru <= 1'b0;
            end
            if(_zz_126) begin
              ways_0_metas_124_mru <= 1'b0;
            end
            if(_zz_127) begin
              ways_0_metas_125_mru <= 1'b0;
            end
            if(_zz_128) begin
              ways_0_metas_126_mru <= 1'b0;
            end
            if(_zz_129) begin
              ways_0_metas_127_mru <= 1'b0;
            end
          end
        end else begin
          if(when_DCache_l224) begin
            if(_zz_2) begin
              ways_0_metas_0_mru <= 1'b1;
            end
            if(_zz_3) begin
              ways_0_metas_1_mru <= 1'b1;
            end
            if(_zz_4) begin
              ways_0_metas_2_mru <= 1'b1;
            end
            if(_zz_5) begin
              ways_0_metas_3_mru <= 1'b1;
            end
            if(_zz_6) begin
              ways_0_metas_4_mru <= 1'b1;
            end
            if(_zz_7) begin
              ways_0_metas_5_mru <= 1'b1;
            end
            if(_zz_8) begin
              ways_0_metas_6_mru <= 1'b1;
            end
            if(_zz_9) begin
              ways_0_metas_7_mru <= 1'b1;
            end
            if(_zz_10) begin
              ways_0_metas_8_mru <= 1'b1;
            end
            if(_zz_11) begin
              ways_0_metas_9_mru <= 1'b1;
            end
            if(_zz_12) begin
              ways_0_metas_10_mru <= 1'b1;
            end
            if(_zz_13) begin
              ways_0_metas_11_mru <= 1'b1;
            end
            if(_zz_14) begin
              ways_0_metas_12_mru <= 1'b1;
            end
            if(_zz_15) begin
              ways_0_metas_13_mru <= 1'b1;
            end
            if(_zz_16) begin
              ways_0_metas_14_mru <= 1'b1;
            end
            if(_zz_17) begin
              ways_0_metas_15_mru <= 1'b1;
            end
            if(_zz_18) begin
              ways_0_metas_16_mru <= 1'b1;
            end
            if(_zz_19) begin
              ways_0_metas_17_mru <= 1'b1;
            end
            if(_zz_20) begin
              ways_0_metas_18_mru <= 1'b1;
            end
            if(_zz_21) begin
              ways_0_metas_19_mru <= 1'b1;
            end
            if(_zz_22) begin
              ways_0_metas_20_mru <= 1'b1;
            end
            if(_zz_23) begin
              ways_0_metas_21_mru <= 1'b1;
            end
            if(_zz_24) begin
              ways_0_metas_22_mru <= 1'b1;
            end
            if(_zz_25) begin
              ways_0_metas_23_mru <= 1'b1;
            end
            if(_zz_26) begin
              ways_0_metas_24_mru <= 1'b1;
            end
            if(_zz_27) begin
              ways_0_metas_25_mru <= 1'b1;
            end
            if(_zz_28) begin
              ways_0_metas_26_mru <= 1'b1;
            end
            if(_zz_29) begin
              ways_0_metas_27_mru <= 1'b1;
            end
            if(_zz_30) begin
              ways_0_metas_28_mru <= 1'b1;
            end
            if(_zz_31) begin
              ways_0_metas_29_mru <= 1'b1;
            end
            if(_zz_32) begin
              ways_0_metas_30_mru <= 1'b1;
            end
            if(_zz_33) begin
              ways_0_metas_31_mru <= 1'b1;
            end
            if(_zz_34) begin
              ways_0_metas_32_mru <= 1'b1;
            end
            if(_zz_35) begin
              ways_0_metas_33_mru <= 1'b1;
            end
            if(_zz_36) begin
              ways_0_metas_34_mru <= 1'b1;
            end
            if(_zz_37) begin
              ways_0_metas_35_mru <= 1'b1;
            end
            if(_zz_38) begin
              ways_0_metas_36_mru <= 1'b1;
            end
            if(_zz_39) begin
              ways_0_metas_37_mru <= 1'b1;
            end
            if(_zz_40) begin
              ways_0_metas_38_mru <= 1'b1;
            end
            if(_zz_41) begin
              ways_0_metas_39_mru <= 1'b1;
            end
            if(_zz_42) begin
              ways_0_metas_40_mru <= 1'b1;
            end
            if(_zz_43) begin
              ways_0_metas_41_mru <= 1'b1;
            end
            if(_zz_44) begin
              ways_0_metas_42_mru <= 1'b1;
            end
            if(_zz_45) begin
              ways_0_metas_43_mru <= 1'b1;
            end
            if(_zz_46) begin
              ways_0_metas_44_mru <= 1'b1;
            end
            if(_zz_47) begin
              ways_0_metas_45_mru <= 1'b1;
            end
            if(_zz_48) begin
              ways_0_metas_46_mru <= 1'b1;
            end
            if(_zz_49) begin
              ways_0_metas_47_mru <= 1'b1;
            end
            if(_zz_50) begin
              ways_0_metas_48_mru <= 1'b1;
            end
            if(_zz_51) begin
              ways_0_metas_49_mru <= 1'b1;
            end
            if(_zz_52) begin
              ways_0_metas_50_mru <= 1'b1;
            end
            if(_zz_53) begin
              ways_0_metas_51_mru <= 1'b1;
            end
            if(_zz_54) begin
              ways_0_metas_52_mru <= 1'b1;
            end
            if(_zz_55) begin
              ways_0_metas_53_mru <= 1'b1;
            end
            if(_zz_56) begin
              ways_0_metas_54_mru <= 1'b1;
            end
            if(_zz_57) begin
              ways_0_metas_55_mru <= 1'b1;
            end
            if(_zz_58) begin
              ways_0_metas_56_mru <= 1'b1;
            end
            if(_zz_59) begin
              ways_0_metas_57_mru <= 1'b1;
            end
            if(_zz_60) begin
              ways_0_metas_58_mru <= 1'b1;
            end
            if(_zz_61) begin
              ways_0_metas_59_mru <= 1'b1;
            end
            if(_zz_62) begin
              ways_0_metas_60_mru <= 1'b1;
            end
            if(_zz_63) begin
              ways_0_metas_61_mru <= 1'b1;
            end
            if(_zz_64) begin
              ways_0_metas_62_mru <= 1'b1;
            end
            if(_zz_65) begin
              ways_0_metas_63_mru <= 1'b1;
            end
            if(_zz_66) begin
              ways_0_metas_64_mru <= 1'b1;
            end
            if(_zz_67) begin
              ways_0_metas_65_mru <= 1'b1;
            end
            if(_zz_68) begin
              ways_0_metas_66_mru <= 1'b1;
            end
            if(_zz_69) begin
              ways_0_metas_67_mru <= 1'b1;
            end
            if(_zz_70) begin
              ways_0_metas_68_mru <= 1'b1;
            end
            if(_zz_71) begin
              ways_0_metas_69_mru <= 1'b1;
            end
            if(_zz_72) begin
              ways_0_metas_70_mru <= 1'b1;
            end
            if(_zz_73) begin
              ways_0_metas_71_mru <= 1'b1;
            end
            if(_zz_74) begin
              ways_0_metas_72_mru <= 1'b1;
            end
            if(_zz_75) begin
              ways_0_metas_73_mru <= 1'b1;
            end
            if(_zz_76) begin
              ways_0_metas_74_mru <= 1'b1;
            end
            if(_zz_77) begin
              ways_0_metas_75_mru <= 1'b1;
            end
            if(_zz_78) begin
              ways_0_metas_76_mru <= 1'b1;
            end
            if(_zz_79) begin
              ways_0_metas_77_mru <= 1'b1;
            end
            if(_zz_80) begin
              ways_0_metas_78_mru <= 1'b1;
            end
            if(_zz_81) begin
              ways_0_metas_79_mru <= 1'b1;
            end
            if(_zz_82) begin
              ways_0_metas_80_mru <= 1'b1;
            end
            if(_zz_83) begin
              ways_0_metas_81_mru <= 1'b1;
            end
            if(_zz_84) begin
              ways_0_metas_82_mru <= 1'b1;
            end
            if(_zz_85) begin
              ways_0_metas_83_mru <= 1'b1;
            end
            if(_zz_86) begin
              ways_0_metas_84_mru <= 1'b1;
            end
            if(_zz_87) begin
              ways_0_metas_85_mru <= 1'b1;
            end
            if(_zz_88) begin
              ways_0_metas_86_mru <= 1'b1;
            end
            if(_zz_89) begin
              ways_0_metas_87_mru <= 1'b1;
            end
            if(_zz_90) begin
              ways_0_metas_88_mru <= 1'b1;
            end
            if(_zz_91) begin
              ways_0_metas_89_mru <= 1'b1;
            end
            if(_zz_92) begin
              ways_0_metas_90_mru <= 1'b1;
            end
            if(_zz_93) begin
              ways_0_metas_91_mru <= 1'b1;
            end
            if(_zz_94) begin
              ways_0_metas_92_mru <= 1'b1;
            end
            if(_zz_95) begin
              ways_0_metas_93_mru <= 1'b1;
            end
            if(_zz_96) begin
              ways_0_metas_94_mru <= 1'b1;
            end
            if(_zz_97) begin
              ways_0_metas_95_mru <= 1'b1;
            end
            if(_zz_98) begin
              ways_0_metas_96_mru <= 1'b1;
            end
            if(_zz_99) begin
              ways_0_metas_97_mru <= 1'b1;
            end
            if(_zz_100) begin
              ways_0_metas_98_mru <= 1'b1;
            end
            if(_zz_101) begin
              ways_0_metas_99_mru <= 1'b1;
            end
            if(_zz_102) begin
              ways_0_metas_100_mru <= 1'b1;
            end
            if(_zz_103) begin
              ways_0_metas_101_mru <= 1'b1;
            end
            if(_zz_104) begin
              ways_0_metas_102_mru <= 1'b1;
            end
            if(_zz_105) begin
              ways_0_metas_103_mru <= 1'b1;
            end
            if(_zz_106) begin
              ways_0_metas_104_mru <= 1'b1;
            end
            if(_zz_107) begin
              ways_0_metas_105_mru <= 1'b1;
            end
            if(_zz_108) begin
              ways_0_metas_106_mru <= 1'b1;
            end
            if(_zz_109) begin
              ways_0_metas_107_mru <= 1'b1;
            end
            if(_zz_110) begin
              ways_0_metas_108_mru <= 1'b1;
            end
            if(_zz_111) begin
              ways_0_metas_109_mru <= 1'b1;
            end
            if(_zz_112) begin
              ways_0_metas_110_mru <= 1'b1;
            end
            if(_zz_113) begin
              ways_0_metas_111_mru <= 1'b1;
            end
            if(_zz_114) begin
              ways_0_metas_112_mru <= 1'b1;
            end
            if(_zz_115) begin
              ways_0_metas_113_mru <= 1'b1;
            end
            if(_zz_116) begin
              ways_0_metas_114_mru <= 1'b1;
            end
            if(_zz_117) begin
              ways_0_metas_115_mru <= 1'b1;
            end
            if(_zz_118) begin
              ways_0_metas_116_mru <= 1'b1;
            end
            if(_zz_119) begin
              ways_0_metas_117_mru <= 1'b1;
            end
            if(_zz_120) begin
              ways_0_metas_118_mru <= 1'b1;
            end
            if(_zz_121) begin
              ways_0_metas_119_mru <= 1'b1;
            end
            if(_zz_122) begin
              ways_0_metas_120_mru <= 1'b1;
            end
            if(_zz_123) begin
              ways_0_metas_121_mru <= 1'b1;
            end
            if(_zz_124) begin
              ways_0_metas_122_mru <= 1'b1;
            end
            if(_zz_125) begin
              ways_0_metas_123_mru <= 1'b1;
            end
            if(_zz_126) begin
              ways_0_metas_124_mru <= 1'b1;
            end
            if(_zz_127) begin
              ways_0_metas_125_mru <= 1'b1;
            end
            if(_zz_128) begin
              ways_0_metas_126_mru <= 1'b1;
            end
            if(_zz_129) begin
              ways_0_metas_127_mru <= 1'b1;
            end
          end else begin
            if(when_DCache_l227) begin
              if(_zz_2) begin
                ways_0_metas_0_vld <= 1'b1;
              end
              if(_zz_3) begin
                ways_0_metas_1_vld <= 1'b1;
              end
              if(_zz_4) begin
                ways_0_metas_2_vld <= 1'b1;
              end
              if(_zz_5) begin
                ways_0_metas_3_vld <= 1'b1;
              end
              if(_zz_6) begin
                ways_0_metas_4_vld <= 1'b1;
              end
              if(_zz_7) begin
                ways_0_metas_5_vld <= 1'b1;
              end
              if(_zz_8) begin
                ways_0_metas_6_vld <= 1'b1;
              end
              if(_zz_9) begin
                ways_0_metas_7_vld <= 1'b1;
              end
              if(_zz_10) begin
                ways_0_metas_8_vld <= 1'b1;
              end
              if(_zz_11) begin
                ways_0_metas_9_vld <= 1'b1;
              end
              if(_zz_12) begin
                ways_0_metas_10_vld <= 1'b1;
              end
              if(_zz_13) begin
                ways_0_metas_11_vld <= 1'b1;
              end
              if(_zz_14) begin
                ways_0_metas_12_vld <= 1'b1;
              end
              if(_zz_15) begin
                ways_0_metas_13_vld <= 1'b1;
              end
              if(_zz_16) begin
                ways_0_metas_14_vld <= 1'b1;
              end
              if(_zz_17) begin
                ways_0_metas_15_vld <= 1'b1;
              end
              if(_zz_18) begin
                ways_0_metas_16_vld <= 1'b1;
              end
              if(_zz_19) begin
                ways_0_metas_17_vld <= 1'b1;
              end
              if(_zz_20) begin
                ways_0_metas_18_vld <= 1'b1;
              end
              if(_zz_21) begin
                ways_0_metas_19_vld <= 1'b1;
              end
              if(_zz_22) begin
                ways_0_metas_20_vld <= 1'b1;
              end
              if(_zz_23) begin
                ways_0_metas_21_vld <= 1'b1;
              end
              if(_zz_24) begin
                ways_0_metas_22_vld <= 1'b1;
              end
              if(_zz_25) begin
                ways_0_metas_23_vld <= 1'b1;
              end
              if(_zz_26) begin
                ways_0_metas_24_vld <= 1'b1;
              end
              if(_zz_27) begin
                ways_0_metas_25_vld <= 1'b1;
              end
              if(_zz_28) begin
                ways_0_metas_26_vld <= 1'b1;
              end
              if(_zz_29) begin
                ways_0_metas_27_vld <= 1'b1;
              end
              if(_zz_30) begin
                ways_0_metas_28_vld <= 1'b1;
              end
              if(_zz_31) begin
                ways_0_metas_29_vld <= 1'b1;
              end
              if(_zz_32) begin
                ways_0_metas_30_vld <= 1'b1;
              end
              if(_zz_33) begin
                ways_0_metas_31_vld <= 1'b1;
              end
              if(_zz_34) begin
                ways_0_metas_32_vld <= 1'b1;
              end
              if(_zz_35) begin
                ways_0_metas_33_vld <= 1'b1;
              end
              if(_zz_36) begin
                ways_0_metas_34_vld <= 1'b1;
              end
              if(_zz_37) begin
                ways_0_metas_35_vld <= 1'b1;
              end
              if(_zz_38) begin
                ways_0_metas_36_vld <= 1'b1;
              end
              if(_zz_39) begin
                ways_0_metas_37_vld <= 1'b1;
              end
              if(_zz_40) begin
                ways_0_metas_38_vld <= 1'b1;
              end
              if(_zz_41) begin
                ways_0_metas_39_vld <= 1'b1;
              end
              if(_zz_42) begin
                ways_0_metas_40_vld <= 1'b1;
              end
              if(_zz_43) begin
                ways_0_metas_41_vld <= 1'b1;
              end
              if(_zz_44) begin
                ways_0_metas_42_vld <= 1'b1;
              end
              if(_zz_45) begin
                ways_0_metas_43_vld <= 1'b1;
              end
              if(_zz_46) begin
                ways_0_metas_44_vld <= 1'b1;
              end
              if(_zz_47) begin
                ways_0_metas_45_vld <= 1'b1;
              end
              if(_zz_48) begin
                ways_0_metas_46_vld <= 1'b1;
              end
              if(_zz_49) begin
                ways_0_metas_47_vld <= 1'b1;
              end
              if(_zz_50) begin
                ways_0_metas_48_vld <= 1'b1;
              end
              if(_zz_51) begin
                ways_0_metas_49_vld <= 1'b1;
              end
              if(_zz_52) begin
                ways_0_metas_50_vld <= 1'b1;
              end
              if(_zz_53) begin
                ways_0_metas_51_vld <= 1'b1;
              end
              if(_zz_54) begin
                ways_0_metas_52_vld <= 1'b1;
              end
              if(_zz_55) begin
                ways_0_metas_53_vld <= 1'b1;
              end
              if(_zz_56) begin
                ways_0_metas_54_vld <= 1'b1;
              end
              if(_zz_57) begin
                ways_0_metas_55_vld <= 1'b1;
              end
              if(_zz_58) begin
                ways_0_metas_56_vld <= 1'b1;
              end
              if(_zz_59) begin
                ways_0_metas_57_vld <= 1'b1;
              end
              if(_zz_60) begin
                ways_0_metas_58_vld <= 1'b1;
              end
              if(_zz_61) begin
                ways_0_metas_59_vld <= 1'b1;
              end
              if(_zz_62) begin
                ways_0_metas_60_vld <= 1'b1;
              end
              if(_zz_63) begin
                ways_0_metas_61_vld <= 1'b1;
              end
              if(_zz_64) begin
                ways_0_metas_62_vld <= 1'b1;
              end
              if(_zz_65) begin
                ways_0_metas_63_vld <= 1'b1;
              end
              if(_zz_66) begin
                ways_0_metas_64_vld <= 1'b1;
              end
              if(_zz_67) begin
                ways_0_metas_65_vld <= 1'b1;
              end
              if(_zz_68) begin
                ways_0_metas_66_vld <= 1'b1;
              end
              if(_zz_69) begin
                ways_0_metas_67_vld <= 1'b1;
              end
              if(_zz_70) begin
                ways_0_metas_68_vld <= 1'b1;
              end
              if(_zz_71) begin
                ways_0_metas_69_vld <= 1'b1;
              end
              if(_zz_72) begin
                ways_0_metas_70_vld <= 1'b1;
              end
              if(_zz_73) begin
                ways_0_metas_71_vld <= 1'b1;
              end
              if(_zz_74) begin
                ways_0_metas_72_vld <= 1'b1;
              end
              if(_zz_75) begin
                ways_0_metas_73_vld <= 1'b1;
              end
              if(_zz_76) begin
                ways_0_metas_74_vld <= 1'b1;
              end
              if(_zz_77) begin
                ways_0_metas_75_vld <= 1'b1;
              end
              if(_zz_78) begin
                ways_0_metas_76_vld <= 1'b1;
              end
              if(_zz_79) begin
                ways_0_metas_77_vld <= 1'b1;
              end
              if(_zz_80) begin
                ways_0_metas_78_vld <= 1'b1;
              end
              if(_zz_81) begin
                ways_0_metas_79_vld <= 1'b1;
              end
              if(_zz_82) begin
                ways_0_metas_80_vld <= 1'b1;
              end
              if(_zz_83) begin
                ways_0_metas_81_vld <= 1'b1;
              end
              if(_zz_84) begin
                ways_0_metas_82_vld <= 1'b1;
              end
              if(_zz_85) begin
                ways_0_metas_83_vld <= 1'b1;
              end
              if(_zz_86) begin
                ways_0_metas_84_vld <= 1'b1;
              end
              if(_zz_87) begin
                ways_0_metas_85_vld <= 1'b1;
              end
              if(_zz_88) begin
                ways_0_metas_86_vld <= 1'b1;
              end
              if(_zz_89) begin
                ways_0_metas_87_vld <= 1'b1;
              end
              if(_zz_90) begin
                ways_0_metas_88_vld <= 1'b1;
              end
              if(_zz_91) begin
                ways_0_metas_89_vld <= 1'b1;
              end
              if(_zz_92) begin
                ways_0_metas_90_vld <= 1'b1;
              end
              if(_zz_93) begin
                ways_0_metas_91_vld <= 1'b1;
              end
              if(_zz_94) begin
                ways_0_metas_92_vld <= 1'b1;
              end
              if(_zz_95) begin
                ways_0_metas_93_vld <= 1'b1;
              end
              if(_zz_96) begin
                ways_0_metas_94_vld <= 1'b1;
              end
              if(_zz_97) begin
                ways_0_metas_95_vld <= 1'b1;
              end
              if(_zz_98) begin
                ways_0_metas_96_vld <= 1'b1;
              end
              if(_zz_99) begin
                ways_0_metas_97_vld <= 1'b1;
              end
              if(_zz_100) begin
                ways_0_metas_98_vld <= 1'b1;
              end
              if(_zz_101) begin
                ways_0_metas_99_vld <= 1'b1;
              end
              if(_zz_102) begin
                ways_0_metas_100_vld <= 1'b1;
              end
              if(_zz_103) begin
                ways_0_metas_101_vld <= 1'b1;
              end
              if(_zz_104) begin
                ways_0_metas_102_vld <= 1'b1;
              end
              if(_zz_105) begin
                ways_0_metas_103_vld <= 1'b1;
              end
              if(_zz_106) begin
                ways_0_metas_104_vld <= 1'b1;
              end
              if(_zz_107) begin
                ways_0_metas_105_vld <= 1'b1;
              end
              if(_zz_108) begin
                ways_0_metas_106_vld <= 1'b1;
              end
              if(_zz_109) begin
                ways_0_metas_107_vld <= 1'b1;
              end
              if(_zz_110) begin
                ways_0_metas_108_vld <= 1'b1;
              end
              if(_zz_111) begin
                ways_0_metas_109_vld <= 1'b1;
              end
              if(_zz_112) begin
                ways_0_metas_110_vld <= 1'b1;
              end
              if(_zz_113) begin
                ways_0_metas_111_vld <= 1'b1;
              end
              if(_zz_114) begin
                ways_0_metas_112_vld <= 1'b1;
              end
              if(_zz_115) begin
                ways_0_metas_113_vld <= 1'b1;
              end
              if(_zz_116) begin
                ways_0_metas_114_vld <= 1'b1;
              end
              if(_zz_117) begin
                ways_0_metas_115_vld <= 1'b1;
              end
              if(_zz_118) begin
                ways_0_metas_116_vld <= 1'b1;
              end
              if(_zz_119) begin
                ways_0_metas_117_vld <= 1'b1;
              end
              if(_zz_120) begin
                ways_0_metas_118_vld <= 1'b1;
              end
              if(_zz_121) begin
                ways_0_metas_119_vld <= 1'b1;
              end
              if(_zz_122) begin
                ways_0_metas_120_vld <= 1'b1;
              end
              if(_zz_123) begin
                ways_0_metas_121_vld <= 1'b1;
              end
              if(_zz_124) begin
                ways_0_metas_122_vld <= 1'b1;
              end
              if(_zz_125) begin
                ways_0_metas_123_vld <= 1'b1;
              end
              if(_zz_126) begin
                ways_0_metas_124_vld <= 1'b1;
              end
              if(_zz_127) begin
                ways_0_metas_125_vld <= 1'b1;
              end
              if(_zz_128) begin
                ways_0_metas_126_vld <= 1'b1;
              end
              if(_zz_129) begin
                ways_0_metas_127_vld <= 1'b1;
              end
            end
          end
        end
      end
      if(when_DCache_l232) begin
        if(_zz_2) begin
          ways_0_metas_0_tag <= cpu_tag;
        end
        if(_zz_3) begin
          ways_0_metas_1_tag <= cpu_tag;
        end
        if(_zz_4) begin
          ways_0_metas_2_tag <= cpu_tag;
        end
        if(_zz_5) begin
          ways_0_metas_3_tag <= cpu_tag;
        end
        if(_zz_6) begin
          ways_0_metas_4_tag <= cpu_tag;
        end
        if(_zz_7) begin
          ways_0_metas_5_tag <= cpu_tag;
        end
        if(_zz_8) begin
          ways_0_metas_6_tag <= cpu_tag;
        end
        if(_zz_9) begin
          ways_0_metas_7_tag <= cpu_tag;
        end
        if(_zz_10) begin
          ways_0_metas_8_tag <= cpu_tag;
        end
        if(_zz_11) begin
          ways_0_metas_9_tag <= cpu_tag;
        end
        if(_zz_12) begin
          ways_0_metas_10_tag <= cpu_tag;
        end
        if(_zz_13) begin
          ways_0_metas_11_tag <= cpu_tag;
        end
        if(_zz_14) begin
          ways_0_metas_12_tag <= cpu_tag;
        end
        if(_zz_15) begin
          ways_0_metas_13_tag <= cpu_tag;
        end
        if(_zz_16) begin
          ways_0_metas_14_tag <= cpu_tag;
        end
        if(_zz_17) begin
          ways_0_metas_15_tag <= cpu_tag;
        end
        if(_zz_18) begin
          ways_0_metas_16_tag <= cpu_tag;
        end
        if(_zz_19) begin
          ways_0_metas_17_tag <= cpu_tag;
        end
        if(_zz_20) begin
          ways_0_metas_18_tag <= cpu_tag;
        end
        if(_zz_21) begin
          ways_0_metas_19_tag <= cpu_tag;
        end
        if(_zz_22) begin
          ways_0_metas_20_tag <= cpu_tag;
        end
        if(_zz_23) begin
          ways_0_metas_21_tag <= cpu_tag;
        end
        if(_zz_24) begin
          ways_0_metas_22_tag <= cpu_tag;
        end
        if(_zz_25) begin
          ways_0_metas_23_tag <= cpu_tag;
        end
        if(_zz_26) begin
          ways_0_metas_24_tag <= cpu_tag;
        end
        if(_zz_27) begin
          ways_0_metas_25_tag <= cpu_tag;
        end
        if(_zz_28) begin
          ways_0_metas_26_tag <= cpu_tag;
        end
        if(_zz_29) begin
          ways_0_metas_27_tag <= cpu_tag;
        end
        if(_zz_30) begin
          ways_0_metas_28_tag <= cpu_tag;
        end
        if(_zz_31) begin
          ways_0_metas_29_tag <= cpu_tag;
        end
        if(_zz_32) begin
          ways_0_metas_30_tag <= cpu_tag;
        end
        if(_zz_33) begin
          ways_0_metas_31_tag <= cpu_tag;
        end
        if(_zz_34) begin
          ways_0_metas_32_tag <= cpu_tag;
        end
        if(_zz_35) begin
          ways_0_metas_33_tag <= cpu_tag;
        end
        if(_zz_36) begin
          ways_0_metas_34_tag <= cpu_tag;
        end
        if(_zz_37) begin
          ways_0_metas_35_tag <= cpu_tag;
        end
        if(_zz_38) begin
          ways_0_metas_36_tag <= cpu_tag;
        end
        if(_zz_39) begin
          ways_0_metas_37_tag <= cpu_tag;
        end
        if(_zz_40) begin
          ways_0_metas_38_tag <= cpu_tag;
        end
        if(_zz_41) begin
          ways_0_metas_39_tag <= cpu_tag;
        end
        if(_zz_42) begin
          ways_0_metas_40_tag <= cpu_tag;
        end
        if(_zz_43) begin
          ways_0_metas_41_tag <= cpu_tag;
        end
        if(_zz_44) begin
          ways_0_metas_42_tag <= cpu_tag;
        end
        if(_zz_45) begin
          ways_0_metas_43_tag <= cpu_tag;
        end
        if(_zz_46) begin
          ways_0_metas_44_tag <= cpu_tag;
        end
        if(_zz_47) begin
          ways_0_metas_45_tag <= cpu_tag;
        end
        if(_zz_48) begin
          ways_0_metas_46_tag <= cpu_tag;
        end
        if(_zz_49) begin
          ways_0_metas_47_tag <= cpu_tag;
        end
        if(_zz_50) begin
          ways_0_metas_48_tag <= cpu_tag;
        end
        if(_zz_51) begin
          ways_0_metas_49_tag <= cpu_tag;
        end
        if(_zz_52) begin
          ways_0_metas_50_tag <= cpu_tag;
        end
        if(_zz_53) begin
          ways_0_metas_51_tag <= cpu_tag;
        end
        if(_zz_54) begin
          ways_0_metas_52_tag <= cpu_tag;
        end
        if(_zz_55) begin
          ways_0_metas_53_tag <= cpu_tag;
        end
        if(_zz_56) begin
          ways_0_metas_54_tag <= cpu_tag;
        end
        if(_zz_57) begin
          ways_0_metas_55_tag <= cpu_tag;
        end
        if(_zz_58) begin
          ways_0_metas_56_tag <= cpu_tag;
        end
        if(_zz_59) begin
          ways_0_metas_57_tag <= cpu_tag;
        end
        if(_zz_60) begin
          ways_0_metas_58_tag <= cpu_tag;
        end
        if(_zz_61) begin
          ways_0_metas_59_tag <= cpu_tag;
        end
        if(_zz_62) begin
          ways_0_metas_60_tag <= cpu_tag;
        end
        if(_zz_63) begin
          ways_0_metas_61_tag <= cpu_tag;
        end
        if(_zz_64) begin
          ways_0_metas_62_tag <= cpu_tag;
        end
        if(_zz_65) begin
          ways_0_metas_63_tag <= cpu_tag;
        end
        if(_zz_66) begin
          ways_0_metas_64_tag <= cpu_tag;
        end
        if(_zz_67) begin
          ways_0_metas_65_tag <= cpu_tag;
        end
        if(_zz_68) begin
          ways_0_metas_66_tag <= cpu_tag;
        end
        if(_zz_69) begin
          ways_0_metas_67_tag <= cpu_tag;
        end
        if(_zz_70) begin
          ways_0_metas_68_tag <= cpu_tag;
        end
        if(_zz_71) begin
          ways_0_metas_69_tag <= cpu_tag;
        end
        if(_zz_72) begin
          ways_0_metas_70_tag <= cpu_tag;
        end
        if(_zz_73) begin
          ways_0_metas_71_tag <= cpu_tag;
        end
        if(_zz_74) begin
          ways_0_metas_72_tag <= cpu_tag;
        end
        if(_zz_75) begin
          ways_0_metas_73_tag <= cpu_tag;
        end
        if(_zz_76) begin
          ways_0_metas_74_tag <= cpu_tag;
        end
        if(_zz_77) begin
          ways_0_metas_75_tag <= cpu_tag;
        end
        if(_zz_78) begin
          ways_0_metas_76_tag <= cpu_tag;
        end
        if(_zz_79) begin
          ways_0_metas_77_tag <= cpu_tag;
        end
        if(_zz_80) begin
          ways_0_metas_78_tag <= cpu_tag;
        end
        if(_zz_81) begin
          ways_0_metas_79_tag <= cpu_tag;
        end
        if(_zz_82) begin
          ways_0_metas_80_tag <= cpu_tag;
        end
        if(_zz_83) begin
          ways_0_metas_81_tag <= cpu_tag;
        end
        if(_zz_84) begin
          ways_0_metas_82_tag <= cpu_tag;
        end
        if(_zz_85) begin
          ways_0_metas_83_tag <= cpu_tag;
        end
        if(_zz_86) begin
          ways_0_metas_84_tag <= cpu_tag;
        end
        if(_zz_87) begin
          ways_0_metas_85_tag <= cpu_tag;
        end
        if(_zz_88) begin
          ways_0_metas_86_tag <= cpu_tag;
        end
        if(_zz_89) begin
          ways_0_metas_87_tag <= cpu_tag;
        end
        if(_zz_90) begin
          ways_0_metas_88_tag <= cpu_tag;
        end
        if(_zz_91) begin
          ways_0_metas_89_tag <= cpu_tag;
        end
        if(_zz_92) begin
          ways_0_metas_90_tag <= cpu_tag;
        end
        if(_zz_93) begin
          ways_0_metas_91_tag <= cpu_tag;
        end
        if(_zz_94) begin
          ways_0_metas_92_tag <= cpu_tag;
        end
        if(_zz_95) begin
          ways_0_metas_93_tag <= cpu_tag;
        end
        if(_zz_96) begin
          ways_0_metas_94_tag <= cpu_tag;
        end
        if(_zz_97) begin
          ways_0_metas_95_tag <= cpu_tag;
        end
        if(_zz_98) begin
          ways_0_metas_96_tag <= cpu_tag;
        end
        if(_zz_99) begin
          ways_0_metas_97_tag <= cpu_tag;
        end
        if(_zz_100) begin
          ways_0_metas_98_tag <= cpu_tag;
        end
        if(_zz_101) begin
          ways_0_metas_99_tag <= cpu_tag;
        end
        if(_zz_102) begin
          ways_0_metas_100_tag <= cpu_tag;
        end
        if(_zz_103) begin
          ways_0_metas_101_tag <= cpu_tag;
        end
        if(_zz_104) begin
          ways_0_metas_102_tag <= cpu_tag;
        end
        if(_zz_105) begin
          ways_0_metas_103_tag <= cpu_tag;
        end
        if(_zz_106) begin
          ways_0_metas_104_tag <= cpu_tag;
        end
        if(_zz_107) begin
          ways_0_metas_105_tag <= cpu_tag;
        end
        if(_zz_108) begin
          ways_0_metas_106_tag <= cpu_tag;
        end
        if(_zz_109) begin
          ways_0_metas_107_tag <= cpu_tag;
        end
        if(_zz_110) begin
          ways_0_metas_108_tag <= cpu_tag;
        end
        if(_zz_111) begin
          ways_0_metas_109_tag <= cpu_tag;
        end
        if(_zz_112) begin
          ways_0_metas_110_tag <= cpu_tag;
        end
        if(_zz_113) begin
          ways_0_metas_111_tag <= cpu_tag;
        end
        if(_zz_114) begin
          ways_0_metas_112_tag <= cpu_tag;
        end
        if(_zz_115) begin
          ways_0_metas_113_tag <= cpu_tag;
        end
        if(_zz_116) begin
          ways_0_metas_114_tag <= cpu_tag;
        end
        if(_zz_117) begin
          ways_0_metas_115_tag <= cpu_tag;
        end
        if(_zz_118) begin
          ways_0_metas_116_tag <= cpu_tag;
        end
        if(_zz_119) begin
          ways_0_metas_117_tag <= cpu_tag;
        end
        if(_zz_120) begin
          ways_0_metas_118_tag <= cpu_tag;
        end
        if(_zz_121) begin
          ways_0_metas_119_tag <= cpu_tag;
        end
        if(_zz_122) begin
          ways_0_metas_120_tag <= cpu_tag;
        end
        if(_zz_123) begin
          ways_0_metas_121_tag <= cpu_tag;
        end
        if(_zz_124) begin
          ways_0_metas_122_tag <= cpu_tag;
        end
        if(_zz_125) begin
          ways_0_metas_123_tag <= cpu_tag;
        end
        if(_zz_126) begin
          ways_0_metas_124_tag <= cpu_tag;
        end
        if(_zz_127) begin
          ways_0_metas_125_tag <= cpu_tag;
        end
        if(_zz_128) begin
          ways_0_metas_126_tag <= cpu_tag;
        end
        if(_zz_129) begin
          ways_0_metas_127_tag <= cpu_tag;
        end
      end
      if(when_DCache_l237) begin
        cpu_cmd_ready_1 <= 1'b0;
      end else begin
        if(when_DCache_l240) begin
          cpu_cmd_ready_1 <= 1'b1;
        end
      end
      if(flush_busy) begin
        if(_zz_389) begin
          ways_1_metas_0_mru <= 1'b0;
        end
        if(_zz_390) begin
          ways_1_metas_1_mru <= 1'b0;
        end
        if(_zz_391) begin
          ways_1_metas_2_mru <= 1'b0;
        end
        if(_zz_392) begin
          ways_1_metas_3_mru <= 1'b0;
        end
        if(_zz_393) begin
          ways_1_metas_4_mru <= 1'b0;
        end
        if(_zz_394) begin
          ways_1_metas_5_mru <= 1'b0;
        end
        if(_zz_395) begin
          ways_1_metas_6_mru <= 1'b0;
        end
        if(_zz_396) begin
          ways_1_metas_7_mru <= 1'b0;
        end
        if(_zz_397) begin
          ways_1_metas_8_mru <= 1'b0;
        end
        if(_zz_398) begin
          ways_1_metas_9_mru <= 1'b0;
        end
        if(_zz_399) begin
          ways_1_metas_10_mru <= 1'b0;
        end
        if(_zz_400) begin
          ways_1_metas_11_mru <= 1'b0;
        end
        if(_zz_401) begin
          ways_1_metas_12_mru <= 1'b0;
        end
        if(_zz_402) begin
          ways_1_metas_13_mru <= 1'b0;
        end
        if(_zz_403) begin
          ways_1_metas_14_mru <= 1'b0;
        end
        if(_zz_404) begin
          ways_1_metas_15_mru <= 1'b0;
        end
        if(_zz_405) begin
          ways_1_metas_16_mru <= 1'b0;
        end
        if(_zz_406) begin
          ways_1_metas_17_mru <= 1'b0;
        end
        if(_zz_407) begin
          ways_1_metas_18_mru <= 1'b0;
        end
        if(_zz_408) begin
          ways_1_metas_19_mru <= 1'b0;
        end
        if(_zz_409) begin
          ways_1_metas_20_mru <= 1'b0;
        end
        if(_zz_410) begin
          ways_1_metas_21_mru <= 1'b0;
        end
        if(_zz_411) begin
          ways_1_metas_22_mru <= 1'b0;
        end
        if(_zz_412) begin
          ways_1_metas_23_mru <= 1'b0;
        end
        if(_zz_413) begin
          ways_1_metas_24_mru <= 1'b0;
        end
        if(_zz_414) begin
          ways_1_metas_25_mru <= 1'b0;
        end
        if(_zz_415) begin
          ways_1_metas_26_mru <= 1'b0;
        end
        if(_zz_416) begin
          ways_1_metas_27_mru <= 1'b0;
        end
        if(_zz_417) begin
          ways_1_metas_28_mru <= 1'b0;
        end
        if(_zz_418) begin
          ways_1_metas_29_mru <= 1'b0;
        end
        if(_zz_419) begin
          ways_1_metas_30_mru <= 1'b0;
        end
        if(_zz_420) begin
          ways_1_metas_31_mru <= 1'b0;
        end
        if(_zz_421) begin
          ways_1_metas_32_mru <= 1'b0;
        end
        if(_zz_422) begin
          ways_1_metas_33_mru <= 1'b0;
        end
        if(_zz_423) begin
          ways_1_metas_34_mru <= 1'b0;
        end
        if(_zz_424) begin
          ways_1_metas_35_mru <= 1'b0;
        end
        if(_zz_425) begin
          ways_1_metas_36_mru <= 1'b0;
        end
        if(_zz_426) begin
          ways_1_metas_37_mru <= 1'b0;
        end
        if(_zz_427) begin
          ways_1_metas_38_mru <= 1'b0;
        end
        if(_zz_428) begin
          ways_1_metas_39_mru <= 1'b0;
        end
        if(_zz_429) begin
          ways_1_metas_40_mru <= 1'b0;
        end
        if(_zz_430) begin
          ways_1_metas_41_mru <= 1'b0;
        end
        if(_zz_431) begin
          ways_1_metas_42_mru <= 1'b0;
        end
        if(_zz_432) begin
          ways_1_metas_43_mru <= 1'b0;
        end
        if(_zz_433) begin
          ways_1_metas_44_mru <= 1'b0;
        end
        if(_zz_434) begin
          ways_1_metas_45_mru <= 1'b0;
        end
        if(_zz_435) begin
          ways_1_metas_46_mru <= 1'b0;
        end
        if(_zz_436) begin
          ways_1_metas_47_mru <= 1'b0;
        end
        if(_zz_437) begin
          ways_1_metas_48_mru <= 1'b0;
        end
        if(_zz_438) begin
          ways_1_metas_49_mru <= 1'b0;
        end
        if(_zz_439) begin
          ways_1_metas_50_mru <= 1'b0;
        end
        if(_zz_440) begin
          ways_1_metas_51_mru <= 1'b0;
        end
        if(_zz_441) begin
          ways_1_metas_52_mru <= 1'b0;
        end
        if(_zz_442) begin
          ways_1_metas_53_mru <= 1'b0;
        end
        if(_zz_443) begin
          ways_1_metas_54_mru <= 1'b0;
        end
        if(_zz_444) begin
          ways_1_metas_55_mru <= 1'b0;
        end
        if(_zz_445) begin
          ways_1_metas_56_mru <= 1'b0;
        end
        if(_zz_446) begin
          ways_1_metas_57_mru <= 1'b0;
        end
        if(_zz_447) begin
          ways_1_metas_58_mru <= 1'b0;
        end
        if(_zz_448) begin
          ways_1_metas_59_mru <= 1'b0;
        end
        if(_zz_449) begin
          ways_1_metas_60_mru <= 1'b0;
        end
        if(_zz_450) begin
          ways_1_metas_61_mru <= 1'b0;
        end
        if(_zz_451) begin
          ways_1_metas_62_mru <= 1'b0;
        end
        if(_zz_452) begin
          ways_1_metas_63_mru <= 1'b0;
        end
        if(_zz_453) begin
          ways_1_metas_64_mru <= 1'b0;
        end
        if(_zz_454) begin
          ways_1_metas_65_mru <= 1'b0;
        end
        if(_zz_455) begin
          ways_1_metas_66_mru <= 1'b0;
        end
        if(_zz_456) begin
          ways_1_metas_67_mru <= 1'b0;
        end
        if(_zz_457) begin
          ways_1_metas_68_mru <= 1'b0;
        end
        if(_zz_458) begin
          ways_1_metas_69_mru <= 1'b0;
        end
        if(_zz_459) begin
          ways_1_metas_70_mru <= 1'b0;
        end
        if(_zz_460) begin
          ways_1_metas_71_mru <= 1'b0;
        end
        if(_zz_461) begin
          ways_1_metas_72_mru <= 1'b0;
        end
        if(_zz_462) begin
          ways_1_metas_73_mru <= 1'b0;
        end
        if(_zz_463) begin
          ways_1_metas_74_mru <= 1'b0;
        end
        if(_zz_464) begin
          ways_1_metas_75_mru <= 1'b0;
        end
        if(_zz_465) begin
          ways_1_metas_76_mru <= 1'b0;
        end
        if(_zz_466) begin
          ways_1_metas_77_mru <= 1'b0;
        end
        if(_zz_467) begin
          ways_1_metas_78_mru <= 1'b0;
        end
        if(_zz_468) begin
          ways_1_metas_79_mru <= 1'b0;
        end
        if(_zz_469) begin
          ways_1_metas_80_mru <= 1'b0;
        end
        if(_zz_470) begin
          ways_1_metas_81_mru <= 1'b0;
        end
        if(_zz_471) begin
          ways_1_metas_82_mru <= 1'b0;
        end
        if(_zz_472) begin
          ways_1_metas_83_mru <= 1'b0;
        end
        if(_zz_473) begin
          ways_1_metas_84_mru <= 1'b0;
        end
        if(_zz_474) begin
          ways_1_metas_85_mru <= 1'b0;
        end
        if(_zz_475) begin
          ways_1_metas_86_mru <= 1'b0;
        end
        if(_zz_476) begin
          ways_1_metas_87_mru <= 1'b0;
        end
        if(_zz_477) begin
          ways_1_metas_88_mru <= 1'b0;
        end
        if(_zz_478) begin
          ways_1_metas_89_mru <= 1'b0;
        end
        if(_zz_479) begin
          ways_1_metas_90_mru <= 1'b0;
        end
        if(_zz_480) begin
          ways_1_metas_91_mru <= 1'b0;
        end
        if(_zz_481) begin
          ways_1_metas_92_mru <= 1'b0;
        end
        if(_zz_482) begin
          ways_1_metas_93_mru <= 1'b0;
        end
        if(_zz_483) begin
          ways_1_metas_94_mru <= 1'b0;
        end
        if(_zz_484) begin
          ways_1_metas_95_mru <= 1'b0;
        end
        if(_zz_485) begin
          ways_1_metas_96_mru <= 1'b0;
        end
        if(_zz_486) begin
          ways_1_metas_97_mru <= 1'b0;
        end
        if(_zz_487) begin
          ways_1_metas_98_mru <= 1'b0;
        end
        if(_zz_488) begin
          ways_1_metas_99_mru <= 1'b0;
        end
        if(_zz_489) begin
          ways_1_metas_100_mru <= 1'b0;
        end
        if(_zz_490) begin
          ways_1_metas_101_mru <= 1'b0;
        end
        if(_zz_491) begin
          ways_1_metas_102_mru <= 1'b0;
        end
        if(_zz_492) begin
          ways_1_metas_103_mru <= 1'b0;
        end
        if(_zz_493) begin
          ways_1_metas_104_mru <= 1'b0;
        end
        if(_zz_494) begin
          ways_1_metas_105_mru <= 1'b0;
        end
        if(_zz_495) begin
          ways_1_metas_106_mru <= 1'b0;
        end
        if(_zz_496) begin
          ways_1_metas_107_mru <= 1'b0;
        end
        if(_zz_497) begin
          ways_1_metas_108_mru <= 1'b0;
        end
        if(_zz_498) begin
          ways_1_metas_109_mru <= 1'b0;
        end
        if(_zz_499) begin
          ways_1_metas_110_mru <= 1'b0;
        end
        if(_zz_500) begin
          ways_1_metas_111_mru <= 1'b0;
        end
        if(_zz_501) begin
          ways_1_metas_112_mru <= 1'b0;
        end
        if(_zz_502) begin
          ways_1_metas_113_mru <= 1'b0;
        end
        if(_zz_503) begin
          ways_1_metas_114_mru <= 1'b0;
        end
        if(_zz_504) begin
          ways_1_metas_115_mru <= 1'b0;
        end
        if(_zz_505) begin
          ways_1_metas_116_mru <= 1'b0;
        end
        if(_zz_506) begin
          ways_1_metas_117_mru <= 1'b0;
        end
        if(_zz_507) begin
          ways_1_metas_118_mru <= 1'b0;
        end
        if(_zz_508) begin
          ways_1_metas_119_mru <= 1'b0;
        end
        if(_zz_509) begin
          ways_1_metas_120_mru <= 1'b0;
        end
        if(_zz_510) begin
          ways_1_metas_121_mru <= 1'b0;
        end
        if(_zz_511) begin
          ways_1_metas_122_mru <= 1'b0;
        end
        if(_zz_512) begin
          ways_1_metas_123_mru <= 1'b0;
        end
        if(_zz_513) begin
          ways_1_metas_124_mru <= 1'b0;
        end
        if(_zz_514) begin
          ways_1_metas_125_mru <= 1'b0;
        end
        if(_zz_515) begin
          ways_1_metas_126_mru <= 1'b0;
        end
        if(_zz_516) begin
          ways_1_metas_127_mru <= 1'b0;
        end
        if(_zz_389) begin
          ways_1_metas_0_vld <= 1'b0;
        end
        if(_zz_390) begin
          ways_1_metas_1_vld <= 1'b0;
        end
        if(_zz_391) begin
          ways_1_metas_2_vld <= 1'b0;
        end
        if(_zz_392) begin
          ways_1_metas_3_vld <= 1'b0;
        end
        if(_zz_393) begin
          ways_1_metas_4_vld <= 1'b0;
        end
        if(_zz_394) begin
          ways_1_metas_5_vld <= 1'b0;
        end
        if(_zz_395) begin
          ways_1_metas_6_vld <= 1'b0;
        end
        if(_zz_396) begin
          ways_1_metas_7_vld <= 1'b0;
        end
        if(_zz_397) begin
          ways_1_metas_8_vld <= 1'b0;
        end
        if(_zz_398) begin
          ways_1_metas_9_vld <= 1'b0;
        end
        if(_zz_399) begin
          ways_1_metas_10_vld <= 1'b0;
        end
        if(_zz_400) begin
          ways_1_metas_11_vld <= 1'b0;
        end
        if(_zz_401) begin
          ways_1_metas_12_vld <= 1'b0;
        end
        if(_zz_402) begin
          ways_1_metas_13_vld <= 1'b0;
        end
        if(_zz_403) begin
          ways_1_metas_14_vld <= 1'b0;
        end
        if(_zz_404) begin
          ways_1_metas_15_vld <= 1'b0;
        end
        if(_zz_405) begin
          ways_1_metas_16_vld <= 1'b0;
        end
        if(_zz_406) begin
          ways_1_metas_17_vld <= 1'b0;
        end
        if(_zz_407) begin
          ways_1_metas_18_vld <= 1'b0;
        end
        if(_zz_408) begin
          ways_1_metas_19_vld <= 1'b0;
        end
        if(_zz_409) begin
          ways_1_metas_20_vld <= 1'b0;
        end
        if(_zz_410) begin
          ways_1_metas_21_vld <= 1'b0;
        end
        if(_zz_411) begin
          ways_1_metas_22_vld <= 1'b0;
        end
        if(_zz_412) begin
          ways_1_metas_23_vld <= 1'b0;
        end
        if(_zz_413) begin
          ways_1_metas_24_vld <= 1'b0;
        end
        if(_zz_414) begin
          ways_1_metas_25_vld <= 1'b0;
        end
        if(_zz_415) begin
          ways_1_metas_26_vld <= 1'b0;
        end
        if(_zz_416) begin
          ways_1_metas_27_vld <= 1'b0;
        end
        if(_zz_417) begin
          ways_1_metas_28_vld <= 1'b0;
        end
        if(_zz_418) begin
          ways_1_metas_29_vld <= 1'b0;
        end
        if(_zz_419) begin
          ways_1_metas_30_vld <= 1'b0;
        end
        if(_zz_420) begin
          ways_1_metas_31_vld <= 1'b0;
        end
        if(_zz_421) begin
          ways_1_metas_32_vld <= 1'b0;
        end
        if(_zz_422) begin
          ways_1_metas_33_vld <= 1'b0;
        end
        if(_zz_423) begin
          ways_1_metas_34_vld <= 1'b0;
        end
        if(_zz_424) begin
          ways_1_metas_35_vld <= 1'b0;
        end
        if(_zz_425) begin
          ways_1_metas_36_vld <= 1'b0;
        end
        if(_zz_426) begin
          ways_1_metas_37_vld <= 1'b0;
        end
        if(_zz_427) begin
          ways_1_metas_38_vld <= 1'b0;
        end
        if(_zz_428) begin
          ways_1_metas_39_vld <= 1'b0;
        end
        if(_zz_429) begin
          ways_1_metas_40_vld <= 1'b0;
        end
        if(_zz_430) begin
          ways_1_metas_41_vld <= 1'b0;
        end
        if(_zz_431) begin
          ways_1_metas_42_vld <= 1'b0;
        end
        if(_zz_432) begin
          ways_1_metas_43_vld <= 1'b0;
        end
        if(_zz_433) begin
          ways_1_metas_44_vld <= 1'b0;
        end
        if(_zz_434) begin
          ways_1_metas_45_vld <= 1'b0;
        end
        if(_zz_435) begin
          ways_1_metas_46_vld <= 1'b0;
        end
        if(_zz_436) begin
          ways_1_metas_47_vld <= 1'b0;
        end
        if(_zz_437) begin
          ways_1_metas_48_vld <= 1'b0;
        end
        if(_zz_438) begin
          ways_1_metas_49_vld <= 1'b0;
        end
        if(_zz_439) begin
          ways_1_metas_50_vld <= 1'b0;
        end
        if(_zz_440) begin
          ways_1_metas_51_vld <= 1'b0;
        end
        if(_zz_441) begin
          ways_1_metas_52_vld <= 1'b0;
        end
        if(_zz_442) begin
          ways_1_metas_53_vld <= 1'b0;
        end
        if(_zz_443) begin
          ways_1_metas_54_vld <= 1'b0;
        end
        if(_zz_444) begin
          ways_1_metas_55_vld <= 1'b0;
        end
        if(_zz_445) begin
          ways_1_metas_56_vld <= 1'b0;
        end
        if(_zz_446) begin
          ways_1_metas_57_vld <= 1'b0;
        end
        if(_zz_447) begin
          ways_1_metas_58_vld <= 1'b0;
        end
        if(_zz_448) begin
          ways_1_metas_59_vld <= 1'b0;
        end
        if(_zz_449) begin
          ways_1_metas_60_vld <= 1'b0;
        end
        if(_zz_450) begin
          ways_1_metas_61_vld <= 1'b0;
        end
        if(_zz_451) begin
          ways_1_metas_62_vld <= 1'b0;
        end
        if(_zz_452) begin
          ways_1_metas_63_vld <= 1'b0;
        end
        if(_zz_453) begin
          ways_1_metas_64_vld <= 1'b0;
        end
        if(_zz_454) begin
          ways_1_metas_65_vld <= 1'b0;
        end
        if(_zz_455) begin
          ways_1_metas_66_vld <= 1'b0;
        end
        if(_zz_456) begin
          ways_1_metas_67_vld <= 1'b0;
        end
        if(_zz_457) begin
          ways_1_metas_68_vld <= 1'b0;
        end
        if(_zz_458) begin
          ways_1_metas_69_vld <= 1'b0;
        end
        if(_zz_459) begin
          ways_1_metas_70_vld <= 1'b0;
        end
        if(_zz_460) begin
          ways_1_metas_71_vld <= 1'b0;
        end
        if(_zz_461) begin
          ways_1_metas_72_vld <= 1'b0;
        end
        if(_zz_462) begin
          ways_1_metas_73_vld <= 1'b0;
        end
        if(_zz_463) begin
          ways_1_metas_74_vld <= 1'b0;
        end
        if(_zz_464) begin
          ways_1_metas_75_vld <= 1'b0;
        end
        if(_zz_465) begin
          ways_1_metas_76_vld <= 1'b0;
        end
        if(_zz_466) begin
          ways_1_metas_77_vld <= 1'b0;
        end
        if(_zz_467) begin
          ways_1_metas_78_vld <= 1'b0;
        end
        if(_zz_468) begin
          ways_1_metas_79_vld <= 1'b0;
        end
        if(_zz_469) begin
          ways_1_metas_80_vld <= 1'b0;
        end
        if(_zz_470) begin
          ways_1_metas_81_vld <= 1'b0;
        end
        if(_zz_471) begin
          ways_1_metas_82_vld <= 1'b0;
        end
        if(_zz_472) begin
          ways_1_metas_83_vld <= 1'b0;
        end
        if(_zz_473) begin
          ways_1_metas_84_vld <= 1'b0;
        end
        if(_zz_474) begin
          ways_1_metas_85_vld <= 1'b0;
        end
        if(_zz_475) begin
          ways_1_metas_86_vld <= 1'b0;
        end
        if(_zz_476) begin
          ways_1_metas_87_vld <= 1'b0;
        end
        if(_zz_477) begin
          ways_1_metas_88_vld <= 1'b0;
        end
        if(_zz_478) begin
          ways_1_metas_89_vld <= 1'b0;
        end
        if(_zz_479) begin
          ways_1_metas_90_vld <= 1'b0;
        end
        if(_zz_480) begin
          ways_1_metas_91_vld <= 1'b0;
        end
        if(_zz_481) begin
          ways_1_metas_92_vld <= 1'b0;
        end
        if(_zz_482) begin
          ways_1_metas_93_vld <= 1'b0;
        end
        if(_zz_483) begin
          ways_1_metas_94_vld <= 1'b0;
        end
        if(_zz_484) begin
          ways_1_metas_95_vld <= 1'b0;
        end
        if(_zz_485) begin
          ways_1_metas_96_vld <= 1'b0;
        end
        if(_zz_486) begin
          ways_1_metas_97_vld <= 1'b0;
        end
        if(_zz_487) begin
          ways_1_metas_98_vld <= 1'b0;
        end
        if(_zz_488) begin
          ways_1_metas_99_vld <= 1'b0;
        end
        if(_zz_489) begin
          ways_1_metas_100_vld <= 1'b0;
        end
        if(_zz_490) begin
          ways_1_metas_101_vld <= 1'b0;
        end
        if(_zz_491) begin
          ways_1_metas_102_vld <= 1'b0;
        end
        if(_zz_492) begin
          ways_1_metas_103_vld <= 1'b0;
        end
        if(_zz_493) begin
          ways_1_metas_104_vld <= 1'b0;
        end
        if(_zz_494) begin
          ways_1_metas_105_vld <= 1'b0;
        end
        if(_zz_495) begin
          ways_1_metas_106_vld <= 1'b0;
        end
        if(_zz_496) begin
          ways_1_metas_107_vld <= 1'b0;
        end
        if(_zz_497) begin
          ways_1_metas_108_vld <= 1'b0;
        end
        if(_zz_498) begin
          ways_1_metas_109_vld <= 1'b0;
        end
        if(_zz_499) begin
          ways_1_metas_110_vld <= 1'b0;
        end
        if(_zz_500) begin
          ways_1_metas_111_vld <= 1'b0;
        end
        if(_zz_501) begin
          ways_1_metas_112_vld <= 1'b0;
        end
        if(_zz_502) begin
          ways_1_metas_113_vld <= 1'b0;
        end
        if(_zz_503) begin
          ways_1_metas_114_vld <= 1'b0;
        end
        if(_zz_504) begin
          ways_1_metas_115_vld <= 1'b0;
        end
        if(_zz_505) begin
          ways_1_metas_116_vld <= 1'b0;
        end
        if(_zz_506) begin
          ways_1_metas_117_vld <= 1'b0;
        end
        if(_zz_507) begin
          ways_1_metas_118_vld <= 1'b0;
        end
        if(_zz_508) begin
          ways_1_metas_119_vld <= 1'b0;
        end
        if(_zz_509) begin
          ways_1_metas_120_vld <= 1'b0;
        end
        if(_zz_510) begin
          ways_1_metas_121_vld <= 1'b0;
        end
        if(_zz_511) begin
          ways_1_metas_122_vld <= 1'b0;
        end
        if(_zz_512) begin
          ways_1_metas_123_vld <= 1'b0;
        end
        if(_zz_513) begin
          ways_1_metas_124_vld <= 1'b0;
        end
        if(_zz_514) begin
          ways_1_metas_125_vld <= 1'b0;
        end
        if(_zz_515) begin
          ways_1_metas_126_vld <= 1'b0;
        end
        if(_zz_516) begin
          ways_1_metas_127_vld <= 1'b0;
        end
      end else begin
        if(when_DCache_l217_1) begin
          if(cache_hit_1) begin
            if(_zz_260) begin
              ways_1_metas_0_mru <= 1'b1;
            end
            if(_zz_261) begin
              ways_1_metas_1_mru <= 1'b1;
            end
            if(_zz_262) begin
              ways_1_metas_2_mru <= 1'b1;
            end
            if(_zz_263) begin
              ways_1_metas_3_mru <= 1'b1;
            end
            if(_zz_264) begin
              ways_1_metas_4_mru <= 1'b1;
            end
            if(_zz_265) begin
              ways_1_metas_5_mru <= 1'b1;
            end
            if(_zz_266) begin
              ways_1_metas_6_mru <= 1'b1;
            end
            if(_zz_267) begin
              ways_1_metas_7_mru <= 1'b1;
            end
            if(_zz_268) begin
              ways_1_metas_8_mru <= 1'b1;
            end
            if(_zz_269) begin
              ways_1_metas_9_mru <= 1'b1;
            end
            if(_zz_270) begin
              ways_1_metas_10_mru <= 1'b1;
            end
            if(_zz_271) begin
              ways_1_metas_11_mru <= 1'b1;
            end
            if(_zz_272) begin
              ways_1_metas_12_mru <= 1'b1;
            end
            if(_zz_273) begin
              ways_1_metas_13_mru <= 1'b1;
            end
            if(_zz_274) begin
              ways_1_metas_14_mru <= 1'b1;
            end
            if(_zz_275) begin
              ways_1_metas_15_mru <= 1'b1;
            end
            if(_zz_276) begin
              ways_1_metas_16_mru <= 1'b1;
            end
            if(_zz_277) begin
              ways_1_metas_17_mru <= 1'b1;
            end
            if(_zz_278) begin
              ways_1_metas_18_mru <= 1'b1;
            end
            if(_zz_279) begin
              ways_1_metas_19_mru <= 1'b1;
            end
            if(_zz_280) begin
              ways_1_metas_20_mru <= 1'b1;
            end
            if(_zz_281) begin
              ways_1_metas_21_mru <= 1'b1;
            end
            if(_zz_282) begin
              ways_1_metas_22_mru <= 1'b1;
            end
            if(_zz_283) begin
              ways_1_metas_23_mru <= 1'b1;
            end
            if(_zz_284) begin
              ways_1_metas_24_mru <= 1'b1;
            end
            if(_zz_285) begin
              ways_1_metas_25_mru <= 1'b1;
            end
            if(_zz_286) begin
              ways_1_metas_26_mru <= 1'b1;
            end
            if(_zz_287) begin
              ways_1_metas_27_mru <= 1'b1;
            end
            if(_zz_288) begin
              ways_1_metas_28_mru <= 1'b1;
            end
            if(_zz_289) begin
              ways_1_metas_29_mru <= 1'b1;
            end
            if(_zz_290) begin
              ways_1_metas_30_mru <= 1'b1;
            end
            if(_zz_291) begin
              ways_1_metas_31_mru <= 1'b1;
            end
            if(_zz_292) begin
              ways_1_metas_32_mru <= 1'b1;
            end
            if(_zz_293) begin
              ways_1_metas_33_mru <= 1'b1;
            end
            if(_zz_294) begin
              ways_1_metas_34_mru <= 1'b1;
            end
            if(_zz_295) begin
              ways_1_metas_35_mru <= 1'b1;
            end
            if(_zz_296) begin
              ways_1_metas_36_mru <= 1'b1;
            end
            if(_zz_297) begin
              ways_1_metas_37_mru <= 1'b1;
            end
            if(_zz_298) begin
              ways_1_metas_38_mru <= 1'b1;
            end
            if(_zz_299) begin
              ways_1_metas_39_mru <= 1'b1;
            end
            if(_zz_300) begin
              ways_1_metas_40_mru <= 1'b1;
            end
            if(_zz_301) begin
              ways_1_metas_41_mru <= 1'b1;
            end
            if(_zz_302) begin
              ways_1_metas_42_mru <= 1'b1;
            end
            if(_zz_303) begin
              ways_1_metas_43_mru <= 1'b1;
            end
            if(_zz_304) begin
              ways_1_metas_44_mru <= 1'b1;
            end
            if(_zz_305) begin
              ways_1_metas_45_mru <= 1'b1;
            end
            if(_zz_306) begin
              ways_1_metas_46_mru <= 1'b1;
            end
            if(_zz_307) begin
              ways_1_metas_47_mru <= 1'b1;
            end
            if(_zz_308) begin
              ways_1_metas_48_mru <= 1'b1;
            end
            if(_zz_309) begin
              ways_1_metas_49_mru <= 1'b1;
            end
            if(_zz_310) begin
              ways_1_metas_50_mru <= 1'b1;
            end
            if(_zz_311) begin
              ways_1_metas_51_mru <= 1'b1;
            end
            if(_zz_312) begin
              ways_1_metas_52_mru <= 1'b1;
            end
            if(_zz_313) begin
              ways_1_metas_53_mru <= 1'b1;
            end
            if(_zz_314) begin
              ways_1_metas_54_mru <= 1'b1;
            end
            if(_zz_315) begin
              ways_1_metas_55_mru <= 1'b1;
            end
            if(_zz_316) begin
              ways_1_metas_56_mru <= 1'b1;
            end
            if(_zz_317) begin
              ways_1_metas_57_mru <= 1'b1;
            end
            if(_zz_318) begin
              ways_1_metas_58_mru <= 1'b1;
            end
            if(_zz_319) begin
              ways_1_metas_59_mru <= 1'b1;
            end
            if(_zz_320) begin
              ways_1_metas_60_mru <= 1'b1;
            end
            if(_zz_321) begin
              ways_1_metas_61_mru <= 1'b1;
            end
            if(_zz_322) begin
              ways_1_metas_62_mru <= 1'b1;
            end
            if(_zz_323) begin
              ways_1_metas_63_mru <= 1'b1;
            end
            if(_zz_324) begin
              ways_1_metas_64_mru <= 1'b1;
            end
            if(_zz_325) begin
              ways_1_metas_65_mru <= 1'b1;
            end
            if(_zz_326) begin
              ways_1_metas_66_mru <= 1'b1;
            end
            if(_zz_327) begin
              ways_1_metas_67_mru <= 1'b1;
            end
            if(_zz_328) begin
              ways_1_metas_68_mru <= 1'b1;
            end
            if(_zz_329) begin
              ways_1_metas_69_mru <= 1'b1;
            end
            if(_zz_330) begin
              ways_1_metas_70_mru <= 1'b1;
            end
            if(_zz_331) begin
              ways_1_metas_71_mru <= 1'b1;
            end
            if(_zz_332) begin
              ways_1_metas_72_mru <= 1'b1;
            end
            if(_zz_333) begin
              ways_1_metas_73_mru <= 1'b1;
            end
            if(_zz_334) begin
              ways_1_metas_74_mru <= 1'b1;
            end
            if(_zz_335) begin
              ways_1_metas_75_mru <= 1'b1;
            end
            if(_zz_336) begin
              ways_1_metas_76_mru <= 1'b1;
            end
            if(_zz_337) begin
              ways_1_metas_77_mru <= 1'b1;
            end
            if(_zz_338) begin
              ways_1_metas_78_mru <= 1'b1;
            end
            if(_zz_339) begin
              ways_1_metas_79_mru <= 1'b1;
            end
            if(_zz_340) begin
              ways_1_metas_80_mru <= 1'b1;
            end
            if(_zz_341) begin
              ways_1_metas_81_mru <= 1'b1;
            end
            if(_zz_342) begin
              ways_1_metas_82_mru <= 1'b1;
            end
            if(_zz_343) begin
              ways_1_metas_83_mru <= 1'b1;
            end
            if(_zz_344) begin
              ways_1_metas_84_mru <= 1'b1;
            end
            if(_zz_345) begin
              ways_1_metas_85_mru <= 1'b1;
            end
            if(_zz_346) begin
              ways_1_metas_86_mru <= 1'b1;
            end
            if(_zz_347) begin
              ways_1_metas_87_mru <= 1'b1;
            end
            if(_zz_348) begin
              ways_1_metas_88_mru <= 1'b1;
            end
            if(_zz_349) begin
              ways_1_metas_89_mru <= 1'b1;
            end
            if(_zz_350) begin
              ways_1_metas_90_mru <= 1'b1;
            end
            if(_zz_351) begin
              ways_1_metas_91_mru <= 1'b1;
            end
            if(_zz_352) begin
              ways_1_metas_92_mru <= 1'b1;
            end
            if(_zz_353) begin
              ways_1_metas_93_mru <= 1'b1;
            end
            if(_zz_354) begin
              ways_1_metas_94_mru <= 1'b1;
            end
            if(_zz_355) begin
              ways_1_metas_95_mru <= 1'b1;
            end
            if(_zz_356) begin
              ways_1_metas_96_mru <= 1'b1;
            end
            if(_zz_357) begin
              ways_1_metas_97_mru <= 1'b1;
            end
            if(_zz_358) begin
              ways_1_metas_98_mru <= 1'b1;
            end
            if(_zz_359) begin
              ways_1_metas_99_mru <= 1'b1;
            end
            if(_zz_360) begin
              ways_1_metas_100_mru <= 1'b1;
            end
            if(_zz_361) begin
              ways_1_metas_101_mru <= 1'b1;
            end
            if(_zz_362) begin
              ways_1_metas_102_mru <= 1'b1;
            end
            if(_zz_363) begin
              ways_1_metas_103_mru <= 1'b1;
            end
            if(_zz_364) begin
              ways_1_metas_104_mru <= 1'b1;
            end
            if(_zz_365) begin
              ways_1_metas_105_mru <= 1'b1;
            end
            if(_zz_366) begin
              ways_1_metas_106_mru <= 1'b1;
            end
            if(_zz_367) begin
              ways_1_metas_107_mru <= 1'b1;
            end
            if(_zz_368) begin
              ways_1_metas_108_mru <= 1'b1;
            end
            if(_zz_369) begin
              ways_1_metas_109_mru <= 1'b1;
            end
            if(_zz_370) begin
              ways_1_metas_110_mru <= 1'b1;
            end
            if(_zz_371) begin
              ways_1_metas_111_mru <= 1'b1;
            end
            if(_zz_372) begin
              ways_1_metas_112_mru <= 1'b1;
            end
            if(_zz_373) begin
              ways_1_metas_113_mru <= 1'b1;
            end
            if(_zz_374) begin
              ways_1_metas_114_mru <= 1'b1;
            end
            if(_zz_375) begin
              ways_1_metas_115_mru <= 1'b1;
            end
            if(_zz_376) begin
              ways_1_metas_116_mru <= 1'b1;
            end
            if(_zz_377) begin
              ways_1_metas_117_mru <= 1'b1;
            end
            if(_zz_378) begin
              ways_1_metas_118_mru <= 1'b1;
            end
            if(_zz_379) begin
              ways_1_metas_119_mru <= 1'b1;
            end
            if(_zz_380) begin
              ways_1_metas_120_mru <= 1'b1;
            end
            if(_zz_381) begin
              ways_1_metas_121_mru <= 1'b1;
            end
            if(_zz_382) begin
              ways_1_metas_122_mru <= 1'b1;
            end
            if(_zz_383) begin
              ways_1_metas_123_mru <= 1'b1;
            end
            if(_zz_384) begin
              ways_1_metas_124_mru <= 1'b1;
            end
            if(_zz_385) begin
              ways_1_metas_125_mru <= 1'b1;
            end
            if(_zz_386) begin
              ways_1_metas_126_mru <= 1'b1;
            end
            if(_zz_387) begin
              ways_1_metas_127_mru <= 1'b1;
            end
          end else begin
            if(_zz_260) begin
              ways_1_metas_0_mru <= 1'b0;
            end
            if(_zz_261) begin
              ways_1_metas_1_mru <= 1'b0;
            end
            if(_zz_262) begin
              ways_1_metas_2_mru <= 1'b0;
            end
            if(_zz_263) begin
              ways_1_metas_3_mru <= 1'b0;
            end
            if(_zz_264) begin
              ways_1_metas_4_mru <= 1'b0;
            end
            if(_zz_265) begin
              ways_1_metas_5_mru <= 1'b0;
            end
            if(_zz_266) begin
              ways_1_metas_6_mru <= 1'b0;
            end
            if(_zz_267) begin
              ways_1_metas_7_mru <= 1'b0;
            end
            if(_zz_268) begin
              ways_1_metas_8_mru <= 1'b0;
            end
            if(_zz_269) begin
              ways_1_metas_9_mru <= 1'b0;
            end
            if(_zz_270) begin
              ways_1_metas_10_mru <= 1'b0;
            end
            if(_zz_271) begin
              ways_1_metas_11_mru <= 1'b0;
            end
            if(_zz_272) begin
              ways_1_metas_12_mru <= 1'b0;
            end
            if(_zz_273) begin
              ways_1_metas_13_mru <= 1'b0;
            end
            if(_zz_274) begin
              ways_1_metas_14_mru <= 1'b0;
            end
            if(_zz_275) begin
              ways_1_metas_15_mru <= 1'b0;
            end
            if(_zz_276) begin
              ways_1_metas_16_mru <= 1'b0;
            end
            if(_zz_277) begin
              ways_1_metas_17_mru <= 1'b0;
            end
            if(_zz_278) begin
              ways_1_metas_18_mru <= 1'b0;
            end
            if(_zz_279) begin
              ways_1_metas_19_mru <= 1'b0;
            end
            if(_zz_280) begin
              ways_1_metas_20_mru <= 1'b0;
            end
            if(_zz_281) begin
              ways_1_metas_21_mru <= 1'b0;
            end
            if(_zz_282) begin
              ways_1_metas_22_mru <= 1'b0;
            end
            if(_zz_283) begin
              ways_1_metas_23_mru <= 1'b0;
            end
            if(_zz_284) begin
              ways_1_metas_24_mru <= 1'b0;
            end
            if(_zz_285) begin
              ways_1_metas_25_mru <= 1'b0;
            end
            if(_zz_286) begin
              ways_1_metas_26_mru <= 1'b0;
            end
            if(_zz_287) begin
              ways_1_metas_27_mru <= 1'b0;
            end
            if(_zz_288) begin
              ways_1_metas_28_mru <= 1'b0;
            end
            if(_zz_289) begin
              ways_1_metas_29_mru <= 1'b0;
            end
            if(_zz_290) begin
              ways_1_metas_30_mru <= 1'b0;
            end
            if(_zz_291) begin
              ways_1_metas_31_mru <= 1'b0;
            end
            if(_zz_292) begin
              ways_1_metas_32_mru <= 1'b0;
            end
            if(_zz_293) begin
              ways_1_metas_33_mru <= 1'b0;
            end
            if(_zz_294) begin
              ways_1_metas_34_mru <= 1'b0;
            end
            if(_zz_295) begin
              ways_1_metas_35_mru <= 1'b0;
            end
            if(_zz_296) begin
              ways_1_metas_36_mru <= 1'b0;
            end
            if(_zz_297) begin
              ways_1_metas_37_mru <= 1'b0;
            end
            if(_zz_298) begin
              ways_1_metas_38_mru <= 1'b0;
            end
            if(_zz_299) begin
              ways_1_metas_39_mru <= 1'b0;
            end
            if(_zz_300) begin
              ways_1_metas_40_mru <= 1'b0;
            end
            if(_zz_301) begin
              ways_1_metas_41_mru <= 1'b0;
            end
            if(_zz_302) begin
              ways_1_metas_42_mru <= 1'b0;
            end
            if(_zz_303) begin
              ways_1_metas_43_mru <= 1'b0;
            end
            if(_zz_304) begin
              ways_1_metas_44_mru <= 1'b0;
            end
            if(_zz_305) begin
              ways_1_metas_45_mru <= 1'b0;
            end
            if(_zz_306) begin
              ways_1_metas_46_mru <= 1'b0;
            end
            if(_zz_307) begin
              ways_1_metas_47_mru <= 1'b0;
            end
            if(_zz_308) begin
              ways_1_metas_48_mru <= 1'b0;
            end
            if(_zz_309) begin
              ways_1_metas_49_mru <= 1'b0;
            end
            if(_zz_310) begin
              ways_1_metas_50_mru <= 1'b0;
            end
            if(_zz_311) begin
              ways_1_metas_51_mru <= 1'b0;
            end
            if(_zz_312) begin
              ways_1_metas_52_mru <= 1'b0;
            end
            if(_zz_313) begin
              ways_1_metas_53_mru <= 1'b0;
            end
            if(_zz_314) begin
              ways_1_metas_54_mru <= 1'b0;
            end
            if(_zz_315) begin
              ways_1_metas_55_mru <= 1'b0;
            end
            if(_zz_316) begin
              ways_1_metas_56_mru <= 1'b0;
            end
            if(_zz_317) begin
              ways_1_metas_57_mru <= 1'b0;
            end
            if(_zz_318) begin
              ways_1_metas_58_mru <= 1'b0;
            end
            if(_zz_319) begin
              ways_1_metas_59_mru <= 1'b0;
            end
            if(_zz_320) begin
              ways_1_metas_60_mru <= 1'b0;
            end
            if(_zz_321) begin
              ways_1_metas_61_mru <= 1'b0;
            end
            if(_zz_322) begin
              ways_1_metas_62_mru <= 1'b0;
            end
            if(_zz_323) begin
              ways_1_metas_63_mru <= 1'b0;
            end
            if(_zz_324) begin
              ways_1_metas_64_mru <= 1'b0;
            end
            if(_zz_325) begin
              ways_1_metas_65_mru <= 1'b0;
            end
            if(_zz_326) begin
              ways_1_metas_66_mru <= 1'b0;
            end
            if(_zz_327) begin
              ways_1_metas_67_mru <= 1'b0;
            end
            if(_zz_328) begin
              ways_1_metas_68_mru <= 1'b0;
            end
            if(_zz_329) begin
              ways_1_metas_69_mru <= 1'b0;
            end
            if(_zz_330) begin
              ways_1_metas_70_mru <= 1'b0;
            end
            if(_zz_331) begin
              ways_1_metas_71_mru <= 1'b0;
            end
            if(_zz_332) begin
              ways_1_metas_72_mru <= 1'b0;
            end
            if(_zz_333) begin
              ways_1_metas_73_mru <= 1'b0;
            end
            if(_zz_334) begin
              ways_1_metas_74_mru <= 1'b0;
            end
            if(_zz_335) begin
              ways_1_metas_75_mru <= 1'b0;
            end
            if(_zz_336) begin
              ways_1_metas_76_mru <= 1'b0;
            end
            if(_zz_337) begin
              ways_1_metas_77_mru <= 1'b0;
            end
            if(_zz_338) begin
              ways_1_metas_78_mru <= 1'b0;
            end
            if(_zz_339) begin
              ways_1_metas_79_mru <= 1'b0;
            end
            if(_zz_340) begin
              ways_1_metas_80_mru <= 1'b0;
            end
            if(_zz_341) begin
              ways_1_metas_81_mru <= 1'b0;
            end
            if(_zz_342) begin
              ways_1_metas_82_mru <= 1'b0;
            end
            if(_zz_343) begin
              ways_1_metas_83_mru <= 1'b0;
            end
            if(_zz_344) begin
              ways_1_metas_84_mru <= 1'b0;
            end
            if(_zz_345) begin
              ways_1_metas_85_mru <= 1'b0;
            end
            if(_zz_346) begin
              ways_1_metas_86_mru <= 1'b0;
            end
            if(_zz_347) begin
              ways_1_metas_87_mru <= 1'b0;
            end
            if(_zz_348) begin
              ways_1_metas_88_mru <= 1'b0;
            end
            if(_zz_349) begin
              ways_1_metas_89_mru <= 1'b0;
            end
            if(_zz_350) begin
              ways_1_metas_90_mru <= 1'b0;
            end
            if(_zz_351) begin
              ways_1_metas_91_mru <= 1'b0;
            end
            if(_zz_352) begin
              ways_1_metas_92_mru <= 1'b0;
            end
            if(_zz_353) begin
              ways_1_metas_93_mru <= 1'b0;
            end
            if(_zz_354) begin
              ways_1_metas_94_mru <= 1'b0;
            end
            if(_zz_355) begin
              ways_1_metas_95_mru <= 1'b0;
            end
            if(_zz_356) begin
              ways_1_metas_96_mru <= 1'b0;
            end
            if(_zz_357) begin
              ways_1_metas_97_mru <= 1'b0;
            end
            if(_zz_358) begin
              ways_1_metas_98_mru <= 1'b0;
            end
            if(_zz_359) begin
              ways_1_metas_99_mru <= 1'b0;
            end
            if(_zz_360) begin
              ways_1_metas_100_mru <= 1'b0;
            end
            if(_zz_361) begin
              ways_1_metas_101_mru <= 1'b0;
            end
            if(_zz_362) begin
              ways_1_metas_102_mru <= 1'b0;
            end
            if(_zz_363) begin
              ways_1_metas_103_mru <= 1'b0;
            end
            if(_zz_364) begin
              ways_1_metas_104_mru <= 1'b0;
            end
            if(_zz_365) begin
              ways_1_metas_105_mru <= 1'b0;
            end
            if(_zz_366) begin
              ways_1_metas_106_mru <= 1'b0;
            end
            if(_zz_367) begin
              ways_1_metas_107_mru <= 1'b0;
            end
            if(_zz_368) begin
              ways_1_metas_108_mru <= 1'b0;
            end
            if(_zz_369) begin
              ways_1_metas_109_mru <= 1'b0;
            end
            if(_zz_370) begin
              ways_1_metas_110_mru <= 1'b0;
            end
            if(_zz_371) begin
              ways_1_metas_111_mru <= 1'b0;
            end
            if(_zz_372) begin
              ways_1_metas_112_mru <= 1'b0;
            end
            if(_zz_373) begin
              ways_1_metas_113_mru <= 1'b0;
            end
            if(_zz_374) begin
              ways_1_metas_114_mru <= 1'b0;
            end
            if(_zz_375) begin
              ways_1_metas_115_mru <= 1'b0;
            end
            if(_zz_376) begin
              ways_1_metas_116_mru <= 1'b0;
            end
            if(_zz_377) begin
              ways_1_metas_117_mru <= 1'b0;
            end
            if(_zz_378) begin
              ways_1_metas_118_mru <= 1'b0;
            end
            if(_zz_379) begin
              ways_1_metas_119_mru <= 1'b0;
            end
            if(_zz_380) begin
              ways_1_metas_120_mru <= 1'b0;
            end
            if(_zz_381) begin
              ways_1_metas_121_mru <= 1'b0;
            end
            if(_zz_382) begin
              ways_1_metas_122_mru <= 1'b0;
            end
            if(_zz_383) begin
              ways_1_metas_123_mru <= 1'b0;
            end
            if(_zz_384) begin
              ways_1_metas_124_mru <= 1'b0;
            end
            if(_zz_385) begin
              ways_1_metas_125_mru <= 1'b0;
            end
            if(_zz_386) begin
              ways_1_metas_126_mru <= 1'b0;
            end
            if(_zz_387) begin
              ways_1_metas_127_mru <= 1'b0;
            end
          end
        end else begin
          if(when_DCache_l224_1) begin
            if(_zz_260) begin
              ways_1_metas_0_mru <= 1'b1;
            end
            if(_zz_261) begin
              ways_1_metas_1_mru <= 1'b1;
            end
            if(_zz_262) begin
              ways_1_metas_2_mru <= 1'b1;
            end
            if(_zz_263) begin
              ways_1_metas_3_mru <= 1'b1;
            end
            if(_zz_264) begin
              ways_1_metas_4_mru <= 1'b1;
            end
            if(_zz_265) begin
              ways_1_metas_5_mru <= 1'b1;
            end
            if(_zz_266) begin
              ways_1_metas_6_mru <= 1'b1;
            end
            if(_zz_267) begin
              ways_1_metas_7_mru <= 1'b1;
            end
            if(_zz_268) begin
              ways_1_metas_8_mru <= 1'b1;
            end
            if(_zz_269) begin
              ways_1_metas_9_mru <= 1'b1;
            end
            if(_zz_270) begin
              ways_1_metas_10_mru <= 1'b1;
            end
            if(_zz_271) begin
              ways_1_metas_11_mru <= 1'b1;
            end
            if(_zz_272) begin
              ways_1_metas_12_mru <= 1'b1;
            end
            if(_zz_273) begin
              ways_1_metas_13_mru <= 1'b1;
            end
            if(_zz_274) begin
              ways_1_metas_14_mru <= 1'b1;
            end
            if(_zz_275) begin
              ways_1_metas_15_mru <= 1'b1;
            end
            if(_zz_276) begin
              ways_1_metas_16_mru <= 1'b1;
            end
            if(_zz_277) begin
              ways_1_metas_17_mru <= 1'b1;
            end
            if(_zz_278) begin
              ways_1_metas_18_mru <= 1'b1;
            end
            if(_zz_279) begin
              ways_1_metas_19_mru <= 1'b1;
            end
            if(_zz_280) begin
              ways_1_metas_20_mru <= 1'b1;
            end
            if(_zz_281) begin
              ways_1_metas_21_mru <= 1'b1;
            end
            if(_zz_282) begin
              ways_1_metas_22_mru <= 1'b1;
            end
            if(_zz_283) begin
              ways_1_metas_23_mru <= 1'b1;
            end
            if(_zz_284) begin
              ways_1_metas_24_mru <= 1'b1;
            end
            if(_zz_285) begin
              ways_1_metas_25_mru <= 1'b1;
            end
            if(_zz_286) begin
              ways_1_metas_26_mru <= 1'b1;
            end
            if(_zz_287) begin
              ways_1_metas_27_mru <= 1'b1;
            end
            if(_zz_288) begin
              ways_1_metas_28_mru <= 1'b1;
            end
            if(_zz_289) begin
              ways_1_metas_29_mru <= 1'b1;
            end
            if(_zz_290) begin
              ways_1_metas_30_mru <= 1'b1;
            end
            if(_zz_291) begin
              ways_1_metas_31_mru <= 1'b1;
            end
            if(_zz_292) begin
              ways_1_metas_32_mru <= 1'b1;
            end
            if(_zz_293) begin
              ways_1_metas_33_mru <= 1'b1;
            end
            if(_zz_294) begin
              ways_1_metas_34_mru <= 1'b1;
            end
            if(_zz_295) begin
              ways_1_metas_35_mru <= 1'b1;
            end
            if(_zz_296) begin
              ways_1_metas_36_mru <= 1'b1;
            end
            if(_zz_297) begin
              ways_1_metas_37_mru <= 1'b1;
            end
            if(_zz_298) begin
              ways_1_metas_38_mru <= 1'b1;
            end
            if(_zz_299) begin
              ways_1_metas_39_mru <= 1'b1;
            end
            if(_zz_300) begin
              ways_1_metas_40_mru <= 1'b1;
            end
            if(_zz_301) begin
              ways_1_metas_41_mru <= 1'b1;
            end
            if(_zz_302) begin
              ways_1_metas_42_mru <= 1'b1;
            end
            if(_zz_303) begin
              ways_1_metas_43_mru <= 1'b1;
            end
            if(_zz_304) begin
              ways_1_metas_44_mru <= 1'b1;
            end
            if(_zz_305) begin
              ways_1_metas_45_mru <= 1'b1;
            end
            if(_zz_306) begin
              ways_1_metas_46_mru <= 1'b1;
            end
            if(_zz_307) begin
              ways_1_metas_47_mru <= 1'b1;
            end
            if(_zz_308) begin
              ways_1_metas_48_mru <= 1'b1;
            end
            if(_zz_309) begin
              ways_1_metas_49_mru <= 1'b1;
            end
            if(_zz_310) begin
              ways_1_metas_50_mru <= 1'b1;
            end
            if(_zz_311) begin
              ways_1_metas_51_mru <= 1'b1;
            end
            if(_zz_312) begin
              ways_1_metas_52_mru <= 1'b1;
            end
            if(_zz_313) begin
              ways_1_metas_53_mru <= 1'b1;
            end
            if(_zz_314) begin
              ways_1_metas_54_mru <= 1'b1;
            end
            if(_zz_315) begin
              ways_1_metas_55_mru <= 1'b1;
            end
            if(_zz_316) begin
              ways_1_metas_56_mru <= 1'b1;
            end
            if(_zz_317) begin
              ways_1_metas_57_mru <= 1'b1;
            end
            if(_zz_318) begin
              ways_1_metas_58_mru <= 1'b1;
            end
            if(_zz_319) begin
              ways_1_metas_59_mru <= 1'b1;
            end
            if(_zz_320) begin
              ways_1_metas_60_mru <= 1'b1;
            end
            if(_zz_321) begin
              ways_1_metas_61_mru <= 1'b1;
            end
            if(_zz_322) begin
              ways_1_metas_62_mru <= 1'b1;
            end
            if(_zz_323) begin
              ways_1_metas_63_mru <= 1'b1;
            end
            if(_zz_324) begin
              ways_1_metas_64_mru <= 1'b1;
            end
            if(_zz_325) begin
              ways_1_metas_65_mru <= 1'b1;
            end
            if(_zz_326) begin
              ways_1_metas_66_mru <= 1'b1;
            end
            if(_zz_327) begin
              ways_1_metas_67_mru <= 1'b1;
            end
            if(_zz_328) begin
              ways_1_metas_68_mru <= 1'b1;
            end
            if(_zz_329) begin
              ways_1_metas_69_mru <= 1'b1;
            end
            if(_zz_330) begin
              ways_1_metas_70_mru <= 1'b1;
            end
            if(_zz_331) begin
              ways_1_metas_71_mru <= 1'b1;
            end
            if(_zz_332) begin
              ways_1_metas_72_mru <= 1'b1;
            end
            if(_zz_333) begin
              ways_1_metas_73_mru <= 1'b1;
            end
            if(_zz_334) begin
              ways_1_metas_74_mru <= 1'b1;
            end
            if(_zz_335) begin
              ways_1_metas_75_mru <= 1'b1;
            end
            if(_zz_336) begin
              ways_1_metas_76_mru <= 1'b1;
            end
            if(_zz_337) begin
              ways_1_metas_77_mru <= 1'b1;
            end
            if(_zz_338) begin
              ways_1_metas_78_mru <= 1'b1;
            end
            if(_zz_339) begin
              ways_1_metas_79_mru <= 1'b1;
            end
            if(_zz_340) begin
              ways_1_metas_80_mru <= 1'b1;
            end
            if(_zz_341) begin
              ways_1_metas_81_mru <= 1'b1;
            end
            if(_zz_342) begin
              ways_1_metas_82_mru <= 1'b1;
            end
            if(_zz_343) begin
              ways_1_metas_83_mru <= 1'b1;
            end
            if(_zz_344) begin
              ways_1_metas_84_mru <= 1'b1;
            end
            if(_zz_345) begin
              ways_1_metas_85_mru <= 1'b1;
            end
            if(_zz_346) begin
              ways_1_metas_86_mru <= 1'b1;
            end
            if(_zz_347) begin
              ways_1_metas_87_mru <= 1'b1;
            end
            if(_zz_348) begin
              ways_1_metas_88_mru <= 1'b1;
            end
            if(_zz_349) begin
              ways_1_metas_89_mru <= 1'b1;
            end
            if(_zz_350) begin
              ways_1_metas_90_mru <= 1'b1;
            end
            if(_zz_351) begin
              ways_1_metas_91_mru <= 1'b1;
            end
            if(_zz_352) begin
              ways_1_metas_92_mru <= 1'b1;
            end
            if(_zz_353) begin
              ways_1_metas_93_mru <= 1'b1;
            end
            if(_zz_354) begin
              ways_1_metas_94_mru <= 1'b1;
            end
            if(_zz_355) begin
              ways_1_metas_95_mru <= 1'b1;
            end
            if(_zz_356) begin
              ways_1_metas_96_mru <= 1'b1;
            end
            if(_zz_357) begin
              ways_1_metas_97_mru <= 1'b1;
            end
            if(_zz_358) begin
              ways_1_metas_98_mru <= 1'b1;
            end
            if(_zz_359) begin
              ways_1_metas_99_mru <= 1'b1;
            end
            if(_zz_360) begin
              ways_1_metas_100_mru <= 1'b1;
            end
            if(_zz_361) begin
              ways_1_metas_101_mru <= 1'b1;
            end
            if(_zz_362) begin
              ways_1_metas_102_mru <= 1'b1;
            end
            if(_zz_363) begin
              ways_1_metas_103_mru <= 1'b1;
            end
            if(_zz_364) begin
              ways_1_metas_104_mru <= 1'b1;
            end
            if(_zz_365) begin
              ways_1_metas_105_mru <= 1'b1;
            end
            if(_zz_366) begin
              ways_1_metas_106_mru <= 1'b1;
            end
            if(_zz_367) begin
              ways_1_metas_107_mru <= 1'b1;
            end
            if(_zz_368) begin
              ways_1_metas_108_mru <= 1'b1;
            end
            if(_zz_369) begin
              ways_1_metas_109_mru <= 1'b1;
            end
            if(_zz_370) begin
              ways_1_metas_110_mru <= 1'b1;
            end
            if(_zz_371) begin
              ways_1_metas_111_mru <= 1'b1;
            end
            if(_zz_372) begin
              ways_1_metas_112_mru <= 1'b1;
            end
            if(_zz_373) begin
              ways_1_metas_113_mru <= 1'b1;
            end
            if(_zz_374) begin
              ways_1_metas_114_mru <= 1'b1;
            end
            if(_zz_375) begin
              ways_1_metas_115_mru <= 1'b1;
            end
            if(_zz_376) begin
              ways_1_metas_116_mru <= 1'b1;
            end
            if(_zz_377) begin
              ways_1_metas_117_mru <= 1'b1;
            end
            if(_zz_378) begin
              ways_1_metas_118_mru <= 1'b1;
            end
            if(_zz_379) begin
              ways_1_metas_119_mru <= 1'b1;
            end
            if(_zz_380) begin
              ways_1_metas_120_mru <= 1'b1;
            end
            if(_zz_381) begin
              ways_1_metas_121_mru <= 1'b1;
            end
            if(_zz_382) begin
              ways_1_metas_122_mru <= 1'b1;
            end
            if(_zz_383) begin
              ways_1_metas_123_mru <= 1'b1;
            end
            if(_zz_384) begin
              ways_1_metas_124_mru <= 1'b1;
            end
            if(_zz_385) begin
              ways_1_metas_125_mru <= 1'b1;
            end
            if(_zz_386) begin
              ways_1_metas_126_mru <= 1'b1;
            end
            if(_zz_387) begin
              ways_1_metas_127_mru <= 1'b1;
            end
          end else begin
            if(when_DCache_l227_1) begin
              if(_zz_260) begin
                ways_1_metas_0_vld <= 1'b1;
              end
              if(_zz_261) begin
                ways_1_metas_1_vld <= 1'b1;
              end
              if(_zz_262) begin
                ways_1_metas_2_vld <= 1'b1;
              end
              if(_zz_263) begin
                ways_1_metas_3_vld <= 1'b1;
              end
              if(_zz_264) begin
                ways_1_metas_4_vld <= 1'b1;
              end
              if(_zz_265) begin
                ways_1_metas_5_vld <= 1'b1;
              end
              if(_zz_266) begin
                ways_1_metas_6_vld <= 1'b1;
              end
              if(_zz_267) begin
                ways_1_metas_7_vld <= 1'b1;
              end
              if(_zz_268) begin
                ways_1_metas_8_vld <= 1'b1;
              end
              if(_zz_269) begin
                ways_1_metas_9_vld <= 1'b1;
              end
              if(_zz_270) begin
                ways_1_metas_10_vld <= 1'b1;
              end
              if(_zz_271) begin
                ways_1_metas_11_vld <= 1'b1;
              end
              if(_zz_272) begin
                ways_1_metas_12_vld <= 1'b1;
              end
              if(_zz_273) begin
                ways_1_metas_13_vld <= 1'b1;
              end
              if(_zz_274) begin
                ways_1_metas_14_vld <= 1'b1;
              end
              if(_zz_275) begin
                ways_1_metas_15_vld <= 1'b1;
              end
              if(_zz_276) begin
                ways_1_metas_16_vld <= 1'b1;
              end
              if(_zz_277) begin
                ways_1_metas_17_vld <= 1'b1;
              end
              if(_zz_278) begin
                ways_1_metas_18_vld <= 1'b1;
              end
              if(_zz_279) begin
                ways_1_metas_19_vld <= 1'b1;
              end
              if(_zz_280) begin
                ways_1_metas_20_vld <= 1'b1;
              end
              if(_zz_281) begin
                ways_1_metas_21_vld <= 1'b1;
              end
              if(_zz_282) begin
                ways_1_metas_22_vld <= 1'b1;
              end
              if(_zz_283) begin
                ways_1_metas_23_vld <= 1'b1;
              end
              if(_zz_284) begin
                ways_1_metas_24_vld <= 1'b1;
              end
              if(_zz_285) begin
                ways_1_metas_25_vld <= 1'b1;
              end
              if(_zz_286) begin
                ways_1_metas_26_vld <= 1'b1;
              end
              if(_zz_287) begin
                ways_1_metas_27_vld <= 1'b1;
              end
              if(_zz_288) begin
                ways_1_metas_28_vld <= 1'b1;
              end
              if(_zz_289) begin
                ways_1_metas_29_vld <= 1'b1;
              end
              if(_zz_290) begin
                ways_1_metas_30_vld <= 1'b1;
              end
              if(_zz_291) begin
                ways_1_metas_31_vld <= 1'b1;
              end
              if(_zz_292) begin
                ways_1_metas_32_vld <= 1'b1;
              end
              if(_zz_293) begin
                ways_1_metas_33_vld <= 1'b1;
              end
              if(_zz_294) begin
                ways_1_metas_34_vld <= 1'b1;
              end
              if(_zz_295) begin
                ways_1_metas_35_vld <= 1'b1;
              end
              if(_zz_296) begin
                ways_1_metas_36_vld <= 1'b1;
              end
              if(_zz_297) begin
                ways_1_metas_37_vld <= 1'b1;
              end
              if(_zz_298) begin
                ways_1_metas_38_vld <= 1'b1;
              end
              if(_zz_299) begin
                ways_1_metas_39_vld <= 1'b1;
              end
              if(_zz_300) begin
                ways_1_metas_40_vld <= 1'b1;
              end
              if(_zz_301) begin
                ways_1_metas_41_vld <= 1'b1;
              end
              if(_zz_302) begin
                ways_1_metas_42_vld <= 1'b1;
              end
              if(_zz_303) begin
                ways_1_metas_43_vld <= 1'b1;
              end
              if(_zz_304) begin
                ways_1_metas_44_vld <= 1'b1;
              end
              if(_zz_305) begin
                ways_1_metas_45_vld <= 1'b1;
              end
              if(_zz_306) begin
                ways_1_metas_46_vld <= 1'b1;
              end
              if(_zz_307) begin
                ways_1_metas_47_vld <= 1'b1;
              end
              if(_zz_308) begin
                ways_1_metas_48_vld <= 1'b1;
              end
              if(_zz_309) begin
                ways_1_metas_49_vld <= 1'b1;
              end
              if(_zz_310) begin
                ways_1_metas_50_vld <= 1'b1;
              end
              if(_zz_311) begin
                ways_1_metas_51_vld <= 1'b1;
              end
              if(_zz_312) begin
                ways_1_metas_52_vld <= 1'b1;
              end
              if(_zz_313) begin
                ways_1_metas_53_vld <= 1'b1;
              end
              if(_zz_314) begin
                ways_1_metas_54_vld <= 1'b1;
              end
              if(_zz_315) begin
                ways_1_metas_55_vld <= 1'b1;
              end
              if(_zz_316) begin
                ways_1_metas_56_vld <= 1'b1;
              end
              if(_zz_317) begin
                ways_1_metas_57_vld <= 1'b1;
              end
              if(_zz_318) begin
                ways_1_metas_58_vld <= 1'b1;
              end
              if(_zz_319) begin
                ways_1_metas_59_vld <= 1'b1;
              end
              if(_zz_320) begin
                ways_1_metas_60_vld <= 1'b1;
              end
              if(_zz_321) begin
                ways_1_metas_61_vld <= 1'b1;
              end
              if(_zz_322) begin
                ways_1_metas_62_vld <= 1'b1;
              end
              if(_zz_323) begin
                ways_1_metas_63_vld <= 1'b1;
              end
              if(_zz_324) begin
                ways_1_metas_64_vld <= 1'b1;
              end
              if(_zz_325) begin
                ways_1_metas_65_vld <= 1'b1;
              end
              if(_zz_326) begin
                ways_1_metas_66_vld <= 1'b1;
              end
              if(_zz_327) begin
                ways_1_metas_67_vld <= 1'b1;
              end
              if(_zz_328) begin
                ways_1_metas_68_vld <= 1'b1;
              end
              if(_zz_329) begin
                ways_1_metas_69_vld <= 1'b1;
              end
              if(_zz_330) begin
                ways_1_metas_70_vld <= 1'b1;
              end
              if(_zz_331) begin
                ways_1_metas_71_vld <= 1'b1;
              end
              if(_zz_332) begin
                ways_1_metas_72_vld <= 1'b1;
              end
              if(_zz_333) begin
                ways_1_metas_73_vld <= 1'b1;
              end
              if(_zz_334) begin
                ways_1_metas_74_vld <= 1'b1;
              end
              if(_zz_335) begin
                ways_1_metas_75_vld <= 1'b1;
              end
              if(_zz_336) begin
                ways_1_metas_76_vld <= 1'b1;
              end
              if(_zz_337) begin
                ways_1_metas_77_vld <= 1'b1;
              end
              if(_zz_338) begin
                ways_1_metas_78_vld <= 1'b1;
              end
              if(_zz_339) begin
                ways_1_metas_79_vld <= 1'b1;
              end
              if(_zz_340) begin
                ways_1_metas_80_vld <= 1'b1;
              end
              if(_zz_341) begin
                ways_1_metas_81_vld <= 1'b1;
              end
              if(_zz_342) begin
                ways_1_metas_82_vld <= 1'b1;
              end
              if(_zz_343) begin
                ways_1_metas_83_vld <= 1'b1;
              end
              if(_zz_344) begin
                ways_1_metas_84_vld <= 1'b1;
              end
              if(_zz_345) begin
                ways_1_metas_85_vld <= 1'b1;
              end
              if(_zz_346) begin
                ways_1_metas_86_vld <= 1'b1;
              end
              if(_zz_347) begin
                ways_1_metas_87_vld <= 1'b1;
              end
              if(_zz_348) begin
                ways_1_metas_88_vld <= 1'b1;
              end
              if(_zz_349) begin
                ways_1_metas_89_vld <= 1'b1;
              end
              if(_zz_350) begin
                ways_1_metas_90_vld <= 1'b1;
              end
              if(_zz_351) begin
                ways_1_metas_91_vld <= 1'b1;
              end
              if(_zz_352) begin
                ways_1_metas_92_vld <= 1'b1;
              end
              if(_zz_353) begin
                ways_1_metas_93_vld <= 1'b1;
              end
              if(_zz_354) begin
                ways_1_metas_94_vld <= 1'b1;
              end
              if(_zz_355) begin
                ways_1_metas_95_vld <= 1'b1;
              end
              if(_zz_356) begin
                ways_1_metas_96_vld <= 1'b1;
              end
              if(_zz_357) begin
                ways_1_metas_97_vld <= 1'b1;
              end
              if(_zz_358) begin
                ways_1_metas_98_vld <= 1'b1;
              end
              if(_zz_359) begin
                ways_1_metas_99_vld <= 1'b1;
              end
              if(_zz_360) begin
                ways_1_metas_100_vld <= 1'b1;
              end
              if(_zz_361) begin
                ways_1_metas_101_vld <= 1'b1;
              end
              if(_zz_362) begin
                ways_1_metas_102_vld <= 1'b1;
              end
              if(_zz_363) begin
                ways_1_metas_103_vld <= 1'b1;
              end
              if(_zz_364) begin
                ways_1_metas_104_vld <= 1'b1;
              end
              if(_zz_365) begin
                ways_1_metas_105_vld <= 1'b1;
              end
              if(_zz_366) begin
                ways_1_metas_106_vld <= 1'b1;
              end
              if(_zz_367) begin
                ways_1_metas_107_vld <= 1'b1;
              end
              if(_zz_368) begin
                ways_1_metas_108_vld <= 1'b1;
              end
              if(_zz_369) begin
                ways_1_metas_109_vld <= 1'b1;
              end
              if(_zz_370) begin
                ways_1_metas_110_vld <= 1'b1;
              end
              if(_zz_371) begin
                ways_1_metas_111_vld <= 1'b1;
              end
              if(_zz_372) begin
                ways_1_metas_112_vld <= 1'b1;
              end
              if(_zz_373) begin
                ways_1_metas_113_vld <= 1'b1;
              end
              if(_zz_374) begin
                ways_1_metas_114_vld <= 1'b1;
              end
              if(_zz_375) begin
                ways_1_metas_115_vld <= 1'b1;
              end
              if(_zz_376) begin
                ways_1_metas_116_vld <= 1'b1;
              end
              if(_zz_377) begin
                ways_1_metas_117_vld <= 1'b1;
              end
              if(_zz_378) begin
                ways_1_metas_118_vld <= 1'b1;
              end
              if(_zz_379) begin
                ways_1_metas_119_vld <= 1'b1;
              end
              if(_zz_380) begin
                ways_1_metas_120_vld <= 1'b1;
              end
              if(_zz_381) begin
                ways_1_metas_121_vld <= 1'b1;
              end
              if(_zz_382) begin
                ways_1_metas_122_vld <= 1'b1;
              end
              if(_zz_383) begin
                ways_1_metas_123_vld <= 1'b1;
              end
              if(_zz_384) begin
                ways_1_metas_124_vld <= 1'b1;
              end
              if(_zz_385) begin
                ways_1_metas_125_vld <= 1'b1;
              end
              if(_zz_386) begin
                ways_1_metas_126_vld <= 1'b1;
              end
              if(_zz_387) begin
                ways_1_metas_127_vld <= 1'b1;
              end
            end
          end
        end
      end
      if(when_DCache_l232_1) begin
        if(_zz_260) begin
          ways_1_metas_0_tag <= cpu_tag;
        end
        if(_zz_261) begin
          ways_1_metas_1_tag <= cpu_tag;
        end
        if(_zz_262) begin
          ways_1_metas_2_tag <= cpu_tag;
        end
        if(_zz_263) begin
          ways_1_metas_3_tag <= cpu_tag;
        end
        if(_zz_264) begin
          ways_1_metas_4_tag <= cpu_tag;
        end
        if(_zz_265) begin
          ways_1_metas_5_tag <= cpu_tag;
        end
        if(_zz_266) begin
          ways_1_metas_6_tag <= cpu_tag;
        end
        if(_zz_267) begin
          ways_1_metas_7_tag <= cpu_tag;
        end
        if(_zz_268) begin
          ways_1_metas_8_tag <= cpu_tag;
        end
        if(_zz_269) begin
          ways_1_metas_9_tag <= cpu_tag;
        end
        if(_zz_270) begin
          ways_1_metas_10_tag <= cpu_tag;
        end
        if(_zz_271) begin
          ways_1_metas_11_tag <= cpu_tag;
        end
        if(_zz_272) begin
          ways_1_metas_12_tag <= cpu_tag;
        end
        if(_zz_273) begin
          ways_1_metas_13_tag <= cpu_tag;
        end
        if(_zz_274) begin
          ways_1_metas_14_tag <= cpu_tag;
        end
        if(_zz_275) begin
          ways_1_metas_15_tag <= cpu_tag;
        end
        if(_zz_276) begin
          ways_1_metas_16_tag <= cpu_tag;
        end
        if(_zz_277) begin
          ways_1_metas_17_tag <= cpu_tag;
        end
        if(_zz_278) begin
          ways_1_metas_18_tag <= cpu_tag;
        end
        if(_zz_279) begin
          ways_1_metas_19_tag <= cpu_tag;
        end
        if(_zz_280) begin
          ways_1_metas_20_tag <= cpu_tag;
        end
        if(_zz_281) begin
          ways_1_metas_21_tag <= cpu_tag;
        end
        if(_zz_282) begin
          ways_1_metas_22_tag <= cpu_tag;
        end
        if(_zz_283) begin
          ways_1_metas_23_tag <= cpu_tag;
        end
        if(_zz_284) begin
          ways_1_metas_24_tag <= cpu_tag;
        end
        if(_zz_285) begin
          ways_1_metas_25_tag <= cpu_tag;
        end
        if(_zz_286) begin
          ways_1_metas_26_tag <= cpu_tag;
        end
        if(_zz_287) begin
          ways_1_metas_27_tag <= cpu_tag;
        end
        if(_zz_288) begin
          ways_1_metas_28_tag <= cpu_tag;
        end
        if(_zz_289) begin
          ways_1_metas_29_tag <= cpu_tag;
        end
        if(_zz_290) begin
          ways_1_metas_30_tag <= cpu_tag;
        end
        if(_zz_291) begin
          ways_1_metas_31_tag <= cpu_tag;
        end
        if(_zz_292) begin
          ways_1_metas_32_tag <= cpu_tag;
        end
        if(_zz_293) begin
          ways_1_metas_33_tag <= cpu_tag;
        end
        if(_zz_294) begin
          ways_1_metas_34_tag <= cpu_tag;
        end
        if(_zz_295) begin
          ways_1_metas_35_tag <= cpu_tag;
        end
        if(_zz_296) begin
          ways_1_metas_36_tag <= cpu_tag;
        end
        if(_zz_297) begin
          ways_1_metas_37_tag <= cpu_tag;
        end
        if(_zz_298) begin
          ways_1_metas_38_tag <= cpu_tag;
        end
        if(_zz_299) begin
          ways_1_metas_39_tag <= cpu_tag;
        end
        if(_zz_300) begin
          ways_1_metas_40_tag <= cpu_tag;
        end
        if(_zz_301) begin
          ways_1_metas_41_tag <= cpu_tag;
        end
        if(_zz_302) begin
          ways_1_metas_42_tag <= cpu_tag;
        end
        if(_zz_303) begin
          ways_1_metas_43_tag <= cpu_tag;
        end
        if(_zz_304) begin
          ways_1_metas_44_tag <= cpu_tag;
        end
        if(_zz_305) begin
          ways_1_metas_45_tag <= cpu_tag;
        end
        if(_zz_306) begin
          ways_1_metas_46_tag <= cpu_tag;
        end
        if(_zz_307) begin
          ways_1_metas_47_tag <= cpu_tag;
        end
        if(_zz_308) begin
          ways_1_metas_48_tag <= cpu_tag;
        end
        if(_zz_309) begin
          ways_1_metas_49_tag <= cpu_tag;
        end
        if(_zz_310) begin
          ways_1_metas_50_tag <= cpu_tag;
        end
        if(_zz_311) begin
          ways_1_metas_51_tag <= cpu_tag;
        end
        if(_zz_312) begin
          ways_1_metas_52_tag <= cpu_tag;
        end
        if(_zz_313) begin
          ways_1_metas_53_tag <= cpu_tag;
        end
        if(_zz_314) begin
          ways_1_metas_54_tag <= cpu_tag;
        end
        if(_zz_315) begin
          ways_1_metas_55_tag <= cpu_tag;
        end
        if(_zz_316) begin
          ways_1_metas_56_tag <= cpu_tag;
        end
        if(_zz_317) begin
          ways_1_metas_57_tag <= cpu_tag;
        end
        if(_zz_318) begin
          ways_1_metas_58_tag <= cpu_tag;
        end
        if(_zz_319) begin
          ways_1_metas_59_tag <= cpu_tag;
        end
        if(_zz_320) begin
          ways_1_metas_60_tag <= cpu_tag;
        end
        if(_zz_321) begin
          ways_1_metas_61_tag <= cpu_tag;
        end
        if(_zz_322) begin
          ways_1_metas_62_tag <= cpu_tag;
        end
        if(_zz_323) begin
          ways_1_metas_63_tag <= cpu_tag;
        end
        if(_zz_324) begin
          ways_1_metas_64_tag <= cpu_tag;
        end
        if(_zz_325) begin
          ways_1_metas_65_tag <= cpu_tag;
        end
        if(_zz_326) begin
          ways_1_metas_66_tag <= cpu_tag;
        end
        if(_zz_327) begin
          ways_1_metas_67_tag <= cpu_tag;
        end
        if(_zz_328) begin
          ways_1_metas_68_tag <= cpu_tag;
        end
        if(_zz_329) begin
          ways_1_metas_69_tag <= cpu_tag;
        end
        if(_zz_330) begin
          ways_1_metas_70_tag <= cpu_tag;
        end
        if(_zz_331) begin
          ways_1_metas_71_tag <= cpu_tag;
        end
        if(_zz_332) begin
          ways_1_metas_72_tag <= cpu_tag;
        end
        if(_zz_333) begin
          ways_1_metas_73_tag <= cpu_tag;
        end
        if(_zz_334) begin
          ways_1_metas_74_tag <= cpu_tag;
        end
        if(_zz_335) begin
          ways_1_metas_75_tag <= cpu_tag;
        end
        if(_zz_336) begin
          ways_1_metas_76_tag <= cpu_tag;
        end
        if(_zz_337) begin
          ways_1_metas_77_tag <= cpu_tag;
        end
        if(_zz_338) begin
          ways_1_metas_78_tag <= cpu_tag;
        end
        if(_zz_339) begin
          ways_1_metas_79_tag <= cpu_tag;
        end
        if(_zz_340) begin
          ways_1_metas_80_tag <= cpu_tag;
        end
        if(_zz_341) begin
          ways_1_metas_81_tag <= cpu_tag;
        end
        if(_zz_342) begin
          ways_1_metas_82_tag <= cpu_tag;
        end
        if(_zz_343) begin
          ways_1_metas_83_tag <= cpu_tag;
        end
        if(_zz_344) begin
          ways_1_metas_84_tag <= cpu_tag;
        end
        if(_zz_345) begin
          ways_1_metas_85_tag <= cpu_tag;
        end
        if(_zz_346) begin
          ways_1_metas_86_tag <= cpu_tag;
        end
        if(_zz_347) begin
          ways_1_metas_87_tag <= cpu_tag;
        end
        if(_zz_348) begin
          ways_1_metas_88_tag <= cpu_tag;
        end
        if(_zz_349) begin
          ways_1_metas_89_tag <= cpu_tag;
        end
        if(_zz_350) begin
          ways_1_metas_90_tag <= cpu_tag;
        end
        if(_zz_351) begin
          ways_1_metas_91_tag <= cpu_tag;
        end
        if(_zz_352) begin
          ways_1_metas_92_tag <= cpu_tag;
        end
        if(_zz_353) begin
          ways_1_metas_93_tag <= cpu_tag;
        end
        if(_zz_354) begin
          ways_1_metas_94_tag <= cpu_tag;
        end
        if(_zz_355) begin
          ways_1_metas_95_tag <= cpu_tag;
        end
        if(_zz_356) begin
          ways_1_metas_96_tag <= cpu_tag;
        end
        if(_zz_357) begin
          ways_1_metas_97_tag <= cpu_tag;
        end
        if(_zz_358) begin
          ways_1_metas_98_tag <= cpu_tag;
        end
        if(_zz_359) begin
          ways_1_metas_99_tag <= cpu_tag;
        end
        if(_zz_360) begin
          ways_1_metas_100_tag <= cpu_tag;
        end
        if(_zz_361) begin
          ways_1_metas_101_tag <= cpu_tag;
        end
        if(_zz_362) begin
          ways_1_metas_102_tag <= cpu_tag;
        end
        if(_zz_363) begin
          ways_1_metas_103_tag <= cpu_tag;
        end
        if(_zz_364) begin
          ways_1_metas_104_tag <= cpu_tag;
        end
        if(_zz_365) begin
          ways_1_metas_105_tag <= cpu_tag;
        end
        if(_zz_366) begin
          ways_1_metas_106_tag <= cpu_tag;
        end
        if(_zz_367) begin
          ways_1_metas_107_tag <= cpu_tag;
        end
        if(_zz_368) begin
          ways_1_metas_108_tag <= cpu_tag;
        end
        if(_zz_369) begin
          ways_1_metas_109_tag <= cpu_tag;
        end
        if(_zz_370) begin
          ways_1_metas_110_tag <= cpu_tag;
        end
        if(_zz_371) begin
          ways_1_metas_111_tag <= cpu_tag;
        end
        if(_zz_372) begin
          ways_1_metas_112_tag <= cpu_tag;
        end
        if(_zz_373) begin
          ways_1_metas_113_tag <= cpu_tag;
        end
        if(_zz_374) begin
          ways_1_metas_114_tag <= cpu_tag;
        end
        if(_zz_375) begin
          ways_1_metas_115_tag <= cpu_tag;
        end
        if(_zz_376) begin
          ways_1_metas_116_tag <= cpu_tag;
        end
        if(_zz_377) begin
          ways_1_metas_117_tag <= cpu_tag;
        end
        if(_zz_378) begin
          ways_1_metas_118_tag <= cpu_tag;
        end
        if(_zz_379) begin
          ways_1_metas_119_tag <= cpu_tag;
        end
        if(_zz_380) begin
          ways_1_metas_120_tag <= cpu_tag;
        end
        if(_zz_381) begin
          ways_1_metas_121_tag <= cpu_tag;
        end
        if(_zz_382) begin
          ways_1_metas_122_tag <= cpu_tag;
        end
        if(_zz_383) begin
          ways_1_metas_123_tag <= cpu_tag;
        end
        if(_zz_384) begin
          ways_1_metas_124_tag <= cpu_tag;
        end
        if(_zz_385) begin
          ways_1_metas_125_tag <= cpu_tag;
        end
        if(_zz_386) begin
          ways_1_metas_126_tag <= cpu_tag;
        end
        if(_zz_387) begin
          ways_1_metas_127_tag <= cpu_tag;
        end
      end
      if(when_DCache_l237_1) begin
        cpu_cmd_ready_1 <= 1'b0;
      end else begin
        if(when_DCache_l240_1) begin
          cpu_cmd_ready_1 <= 1'b1;
        end
      end
      if(flush_busy) begin
        if(_zz_647) begin
          ways_2_metas_0_mru <= 1'b0;
        end
        if(_zz_648) begin
          ways_2_metas_1_mru <= 1'b0;
        end
        if(_zz_649) begin
          ways_2_metas_2_mru <= 1'b0;
        end
        if(_zz_650) begin
          ways_2_metas_3_mru <= 1'b0;
        end
        if(_zz_651) begin
          ways_2_metas_4_mru <= 1'b0;
        end
        if(_zz_652) begin
          ways_2_metas_5_mru <= 1'b0;
        end
        if(_zz_653) begin
          ways_2_metas_6_mru <= 1'b0;
        end
        if(_zz_654) begin
          ways_2_metas_7_mru <= 1'b0;
        end
        if(_zz_655) begin
          ways_2_metas_8_mru <= 1'b0;
        end
        if(_zz_656) begin
          ways_2_metas_9_mru <= 1'b0;
        end
        if(_zz_657) begin
          ways_2_metas_10_mru <= 1'b0;
        end
        if(_zz_658) begin
          ways_2_metas_11_mru <= 1'b0;
        end
        if(_zz_659) begin
          ways_2_metas_12_mru <= 1'b0;
        end
        if(_zz_660) begin
          ways_2_metas_13_mru <= 1'b0;
        end
        if(_zz_661) begin
          ways_2_metas_14_mru <= 1'b0;
        end
        if(_zz_662) begin
          ways_2_metas_15_mru <= 1'b0;
        end
        if(_zz_663) begin
          ways_2_metas_16_mru <= 1'b0;
        end
        if(_zz_664) begin
          ways_2_metas_17_mru <= 1'b0;
        end
        if(_zz_665) begin
          ways_2_metas_18_mru <= 1'b0;
        end
        if(_zz_666) begin
          ways_2_metas_19_mru <= 1'b0;
        end
        if(_zz_667) begin
          ways_2_metas_20_mru <= 1'b0;
        end
        if(_zz_668) begin
          ways_2_metas_21_mru <= 1'b0;
        end
        if(_zz_669) begin
          ways_2_metas_22_mru <= 1'b0;
        end
        if(_zz_670) begin
          ways_2_metas_23_mru <= 1'b0;
        end
        if(_zz_671) begin
          ways_2_metas_24_mru <= 1'b0;
        end
        if(_zz_672) begin
          ways_2_metas_25_mru <= 1'b0;
        end
        if(_zz_673) begin
          ways_2_metas_26_mru <= 1'b0;
        end
        if(_zz_674) begin
          ways_2_metas_27_mru <= 1'b0;
        end
        if(_zz_675) begin
          ways_2_metas_28_mru <= 1'b0;
        end
        if(_zz_676) begin
          ways_2_metas_29_mru <= 1'b0;
        end
        if(_zz_677) begin
          ways_2_metas_30_mru <= 1'b0;
        end
        if(_zz_678) begin
          ways_2_metas_31_mru <= 1'b0;
        end
        if(_zz_679) begin
          ways_2_metas_32_mru <= 1'b0;
        end
        if(_zz_680) begin
          ways_2_metas_33_mru <= 1'b0;
        end
        if(_zz_681) begin
          ways_2_metas_34_mru <= 1'b0;
        end
        if(_zz_682) begin
          ways_2_metas_35_mru <= 1'b0;
        end
        if(_zz_683) begin
          ways_2_metas_36_mru <= 1'b0;
        end
        if(_zz_684) begin
          ways_2_metas_37_mru <= 1'b0;
        end
        if(_zz_685) begin
          ways_2_metas_38_mru <= 1'b0;
        end
        if(_zz_686) begin
          ways_2_metas_39_mru <= 1'b0;
        end
        if(_zz_687) begin
          ways_2_metas_40_mru <= 1'b0;
        end
        if(_zz_688) begin
          ways_2_metas_41_mru <= 1'b0;
        end
        if(_zz_689) begin
          ways_2_metas_42_mru <= 1'b0;
        end
        if(_zz_690) begin
          ways_2_metas_43_mru <= 1'b0;
        end
        if(_zz_691) begin
          ways_2_metas_44_mru <= 1'b0;
        end
        if(_zz_692) begin
          ways_2_metas_45_mru <= 1'b0;
        end
        if(_zz_693) begin
          ways_2_metas_46_mru <= 1'b0;
        end
        if(_zz_694) begin
          ways_2_metas_47_mru <= 1'b0;
        end
        if(_zz_695) begin
          ways_2_metas_48_mru <= 1'b0;
        end
        if(_zz_696) begin
          ways_2_metas_49_mru <= 1'b0;
        end
        if(_zz_697) begin
          ways_2_metas_50_mru <= 1'b0;
        end
        if(_zz_698) begin
          ways_2_metas_51_mru <= 1'b0;
        end
        if(_zz_699) begin
          ways_2_metas_52_mru <= 1'b0;
        end
        if(_zz_700) begin
          ways_2_metas_53_mru <= 1'b0;
        end
        if(_zz_701) begin
          ways_2_metas_54_mru <= 1'b0;
        end
        if(_zz_702) begin
          ways_2_metas_55_mru <= 1'b0;
        end
        if(_zz_703) begin
          ways_2_metas_56_mru <= 1'b0;
        end
        if(_zz_704) begin
          ways_2_metas_57_mru <= 1'b0;
        end
        if(_zz_705) begin
          ways_2_metas_58_mru <= 1'b0;
        end
        if(_zz_706) begin
          ways_2_metas_59_mru <= 1'b0;
        end
        if(_zz_707) begin
          ways_2_metas_60_mru <= 1'b0;
        end
        if(_zz_708) begin
          ways_2_metas_61_mru <= 1'b0;
        end
        if(_zz_709) begin
          ways_2_metas_62_mru <= 1'b0;
        end
        if(_zz_710) begin
          ways_2_metas_63_mru <= 1'b0;
        end
        if(_zz_711) begin
          ways_2_metas_64_mru <= 1'b0;
        end
        if(_zz_712) begin
          ways_2_metas_65_mru <= 1'b0;
        end
        if(_zz_713) begin
          ways_2_metas_66_mru <= 1'b0;
        end
        if(_zz_714) begin
          ways_2_metas_67_mru <= 1'b0;
        end
        if(_zz_715) begin
          ways_2_metas_68_mru <= 1'b0;
        end
        if(_zz_716) begin
          ways_2_metas_69_mru <= 1'b0;
        end
        if(_zz_717) begin
          ways_2_metas_70_mru <= 1'b0;
        end
        if(_zz_718) begin
          ways_2_metas_71_mru <= 1'b0;
        end
        if(_zz_719) begin
          ways_2_metas_72_mru <= 1'b0;
        end
        if(_zz_720) begin
          ways_2_metas_73_mru <= 1'b0;
        end
        if(_zz_721) begin
          ways_2_metas_74_mru <= 1'b0;
        end
        if(_zz_722) begin
          ways_2_metas_75_mru <= 1'b0;
        end
        if(_zz_723) begin
          ways_2_metas_76_mru <= 1'b0;
        end
        if(_zz_724) begin
          ways_2_metas_77_mru <= 1'b0;
        end
        if(_zz_725) begin
          ways_2_metas_78_mru <= 1'b0;
        end
        if(_zz_726) begin
          ways_2_metas_79_mru <= 1'b0;
        end
        if(_zz_727) begin
          ways_2_metas_80_mru <= 1'b0;
        end
        if(_zz_728) begin
          ways_2_metas_81_mru <= 1'b0;
        end
        if(_zz_729) begin
          ways_2_metas_82_mru <= 1'b0;
        end
        if(_zz_730) begin
          ways_2_metas_83_mru <= 1'b0;
        end
        if(_zz_731) begin
          ways_2_metas_84_mru <= 1'b0;
        end
        if(_zz_732) begin
          ways_2_metas_85_mru <= 1'b0;
        end
        if(_zz_733) begin
          ways_2_metas_86_mru <= 1'b0;
        end
        if(_zz_734) begin
          ways_2_metas_87_mru <= 1'b0;
        end
        if(_zz_735) begin
          ways_2_metas_88_mru <= 1'b0;
        end
        if(_zz_736) begin
          ways_2_metas_89_mru <= 1'b0;
        end
        if(_zz_737) begin
          ways_2_metas_90_mru <= 1'b0;
        end
        if(_zz_738) begin
          ways_2_metas_91_mru <= 1'b0;
        end
        if(_zz_739) begin
          ways_2_metas_92_mru <= 1'b0;
        end
        if(_zz_740) begin
          ways_2_metas_93_mru <= 1'b0;
        end
        if(_zz_741) begin
          ways_2_metas_94_mru <= 1'b0;
        end
        if(_zz_742) begin
          ways_2_metas_95_mru <= 1'b0;
        end
        if(_zz_743) begin
          ways_2_metas_96_mru <= 1'b0;
        end
        if(_zz_744) begin
          ways_2_metas_97_mru <= 1'b0;
        end
        if(_zz_745) begin
          ways_2_metas_98_mru <= 1'b0;
        end
        if(_zz_746) begin
          ways_2_metas_99_mru <= 1'b0;
        end
        if(_zz_747) begin
          ways_2_metas_100_mru <= 1'b0;
        end
        if(_zz_748) begin
          ways_2_metas_101_mru <= 1'b0;
        end
        if(_zz_749) begin
          ways_2_metas_102_mru <= 1'b0;
        end
        if(_zz_750) begin
          ways_2_metas_103_mru <= 1'b0;
        end
        if(_zz_751) begin
          ways_2_metas_104_mru <= 1'b0;
        end
        if(_zz_752) begin
          ways_2_metas_105_mru <= 1'b0;
        end
        if(_zz_753) begin
          ways_2_metas_106_mru <= 1'b0;
        end
        if(_zz_754) begin
          ways_2_metas_107_mru <= 1'b0;
        end
        if(_zz_755) begin
          ways_2_metas_108_mru <= 1'b0;
        end
        if(_zz_756) begin
          ways_2_metas_109_mru <= 1'b0;
        end
        if(_zz_757) begin
          ways_2_metas_110_mru <= 1'b0;
        end
        if(_zz_758) begin
          ways_2_metas_111_mru <= 1'b0;
        end
        if(_zz_759) begin
          ways_2_metas_112_mru <= 1'b0;
        end
        if(_zz_760) begin
          ways_2_metas_113_mru <= 1'b0;
        end
        if(_zz_761) begin
          ways_2_metas_114_mru <= 1'b0;
        end
        if(_zz_762) begin
          ways_2_metas_115_mru <= 1'b0;
        end
        if(_zz_763) begin
          ways_2_metas_116_mru <= 1'b0;
        end
        if(_zz_764) begin
          ways_2_metas_117_mru <= 1'b0;
        end
        if(_zz_765) begin
          ways_2_metas_118_mru <= 1'b0;
        end
        if(_zz_766) begin
          ways_2_metas_119_mru <= 1'b0;
        end
        if(_zz_767) begin
          ways_2_metas_120_mru <= 1'b0;
        end
        if(_zz_768) begin
          ways_2_metas_121_mru <= 1'b0;
        end
        if(_zz_769) begin
          ways_2_metas_122_mru <= 1'b0;
        end
        if(_zz_770) begin
          ways_2_metas_123_mru <= 1'b0;
        end
        if(_zz_771) begin
          ways_2_metas_124_mru <= 1'b0;
        end
        if(_zz_772) begin
          ways_2_metas_125_mru <= 1'b0;
        end
        if(_zz_773) begin
          ways_2_metas_126_mru <= 1'b0;
        end
        if(_zz_774) begin
          ways_2_metas_127_mru <= 1'b0;
        end
        if(_zz_647) begin
          ways_2_metas_0_vld <= 1'b0;
        end
        if(_zz_648) begin
          ways_2_metas_1_vld <= 1'b0;
        end
        if(_zz_649) begin
          ways_2_metas_2_vld <= 1'b0;
        end
        if(_zz_650) begin
          ways_2_metas_3_vld <= 1'b0;
        end
        if(_zz_651) begin
          ways_2_metas_4_vld <= 1'b0;
        end
        if(_zz_652) begin
          ways_2_metas_5_vld <= 1'b0;
        end
        if(_zz_653) begin
          ways_2_metas_6_vld <= 1'b0;
        end
        if(_zz_654) begin
          ways_2_metas_7_vld <= 1'b0;
        end
        if(_zz_655) begin
          ways_2_metas_8_vld <= 1'b0;
        end
        if(_zz_656) begin
          ways_2_metas_9_vld <= 1'b0;
        end
        if(_zz_657) begin
          ways_2_metas_10_vld <= 1'b0;
        end
        if(_zz_658) begin
          ways_2_metas_11_vld <= 1'b0;
        end
        if(_zz_659) begin
          ways_2_metas_12_vld <= 1'b0;
        end
        if(_zz_660) begin
          ways_2_metas_13_vld <= 1'b0;
        end
        if(_zz_661) begin
          ways_2_metas_14_vld <= 1'b0;
        end
        if(_zz_662) begin
          ways_2_metas_15_vld <= 1'b0;
        end
        if(_zz_663) begin
          ways_2_metas_16_vld <= 1'b0;
        end
        if(_zz_664) begin
          ways_2_metas_17_vld <= 1'b0;
        end
        if(_zz_665) begin
          ways_2_metas_18_vld <= 1'b0;
        end
        if(_zz_666) begin
          ways_2_metas_19_vld <= 1'b0;
        end
        if(_zz_667) begin
          ways_2_metas_20_vld <= 1'b0;
        end
        if(_zz_668) begin
          ways_2_metas_21_vld <= 1'b0;
        end
        if(_zz_669) begin
          ways_2_metas_22_vld <= 1'b0;
        end
        if(_zz_670) begin
          ways_2_metas_23_vld <= 1'b0;
        end
        if(_zz_671) begin
          ways_2_metas_24_vld <= 1'b0;
        end
        if(_zz_672) begin
          ways_2_metas_25_vld <= 1'b0;
        end
        if(_zz_673) begin
          ways_2_metas_26_vld <= 1'b0;
        end
        if(_zz_674) begin
          ways_2_metas_27_vld <= 1'b0;
        end
        if(_zz_675) begin
          ways_2_metas_28_vld <= 1'b0;
        end
        if(_zz_676) begin
          ways_2_metas_29_vld <= 1'b0;
        end
        if(_zz_677) begin
          ways_2_metas_30_vld <= 1'b0;
        end
        if(_zz_678) begin
          ways_2_metas_31_vld <= 1'b0;
        end
        if(_zz_679) begin
          ways_2_metas_32_vld <= 1'b0;
        end
        if(_zz_680) begin
          ways_2_metas_33_vld <= 1'b0;
        end
        if(_zz_681) begin
          ways_2_metas_34_vld <= 1'b0;
        end
        if(_zz_682) begin
          ways_2_metas_35_vld <= 1'b0;
        end
        if(_zz_683) begin
          ways_2_metas_36_vld <= 1'b0;
        end
        if(_zz_684) begin
          ways_2_metas_37_vld <= 1'b0;
        end
        if(_zz_685) begin
          ways_2_metas_38_vld <= 1'b0;
        end
        if(_zz_686) begin
          ways_2_metas_39_vld <= 1'b0;
        end
        if(_zz_687) begin
          ways_2_metas_40_vld <= 1'b0;
        end
        if(_zz_688) begin
          ways_2_metas_41_vld <= 1'b0;
        end
        if(_zz_689) begin
          ways_2_metas_42_vld <= 1'b0;
        end
        if(_zz_690) begin
          ways_2_metas_43_vld <= 1'b0;
        end
        if(_zz_691) begin
          ways_2_metas_44_vld <= 1'b0;
        end
        if(_zz_692) begin
          ways_2_metas_45_vld <= 1'b0;
        end
        if(_zz_693) begin
          ways_2_metas_46_vld <= 1'b0;
        end
        if(_zz_694) begin
          ways_2_metas_47_vld <= 1'b0;
        end
        if(_zz_695) begin
          ways_2_metas_48_vld <= 1'b0;
        end
        if(_zz_696) begin
          ways_2_metas_49_vld <= 1'b0;
        end
        if(_zz_697) begin
          ways_2_metas_50_vld <= 1'b0;
        end
        if(_zz_698) begin
          ways_2_metas_51_vld <= 1'b0;
        end
        if(_zz_699) begin
          ways_2_metas_52_vld <= 1'b0;
        end
        if(_zz_700) begin
          ways_2_metas_53_vld <= 1'b0;
        end
        if(_zz_701) begin
          ways_2_metas_54_vld <= 1'b0;
        end
        if(_zz_702) begin
          ways_2_metas_55_vld <= 1'b0;
        end
        if(_zz_703) begin
          ways_2_metas_56_vld <= 1'b0;
        end
        if(_zz_704) begin
          ways_2_metas_57_vld <= 1'b0;
        end
        if(_zz_705) begin
          ways_2_metas_58_vld <= 1'b0;
        end
        if(_zz_706) begin
          ways_2_metas_59_vld <= 1'b0;
        end
        if(_zz_707) begin
          ways_2_metas_60_vld <= 1'b0;
        end
        if(_zz_708) begin
          ways_2_metas_61_vld <= 1'b0;
        end
        if(_zz_709) begin
          ways_2_metas_62_vld <= 1'b0;
        end
        if(_zz_710) begin
          ways_2_metas_63_vld <= 1'b0;
        end
        if(_zz_711) begin
          ways_2_metas_64_vld <= 1'b0;
        end
        if(_zz_712) begin
          ways_2_metas_65_vld <= 1'b0;
        end
        if(_zz_713) begin
          ways_2_metas_66_vld <= 1'b0;
        end
        if(_zz_714) begin
          ways_2_metas_67_vld <= 1'b0;
        end
        if(_zz_715) begin
          ways_2_metas_68_vld <= 1'b0;
        end
        if(_zz_716) begin
          ways_2_metas_69_vld <= 1'b0;
        end
        if(_zz_717) begin
          ways_2_metas_70_vld <= 1'b0;
        end
        if(_zz_718) begin
          ways_2_metas_71_vld <= 1'b0;
        end
        if(_zz_719) begin
          ways_2_metas_72_vld <= 1'b0;
        end
        if(_zz_720) begin
          ways_2_metas_73_vld <= 1'b0;
        end
        if(_zz_721) begin
          ways_2_metas_74_vld <= 1'b0;
        end
        if(_zz_722) begin
          ways_2_metas_75_vld <= 1'b0;
        end
        if(_zz_723) begin
          ways_2_metas_76_vld <= 1'b0;
        end
        if(_zz_724) begin
          ways_2_metas_77_vld <= 1'b0;
        end
        if(_zz_725) begin
          ways_2_metas_78_vld <= 1'b0;
        end
        if(_zz_726) begin
          ways_2_metas_79_vld <= 1'b0;
        end
        if(_zz_727) begin
          ways_2_metas_80_vld <= 1'b0;
        end
        if(_zz_728) begin
          ways_2_metas_81_vld <= 1'b0;
        end
        if(_zz_729) begin
          ways_2_metas_82_vld <= 1'b0;
        end
        if(_zz_730) begin
          ways_2_metas_83_vld <= 1'b0;
        end
        if(_zz_731) begin
          ways_2_metas_84_vld <= 1'b0;
        end
        if(_zz_732) begin
          ways_2_metas_85_vld <= 1'b0;
        end
        if(_zz_733) begin
          ways_2_metas_86_vld <= 1'b0;
        end
        if(_zz_734) begin
          ways_2_metas_87_vld <= 1'b0;
        end
        if(_zz_735) begin
          ways_2_metas_88_vld <= 1'b0;
        end
        if(_zz_736) begin
          ways_2_metas_89_vld <= 1'b0;
        end
        if(_zz_737) begin
          ways_2_metas_90_vld <= 1'b0;
        end
        if(_zz_738) begin
          ways_2_metas_91_vld <= 1'b0;
        end
        if(_zz_739) begin
          ways_2_metas_92_vld <= 1'b0;
        end
        if(_zz_740) begin
          ways_2_metas_93_vld <= 1'b0;
        end
        if(_zz_741) begin
          ways_2_metas_94_vld <= 1'b0;
        end
        if(_zz_742) begin
          ways_2_metas_95_vld <= 1'b0;
        end
        if(_zz_743) begin
          ways_2_metas_96_vld <= 1'b0;
        end
        if(_zz_744) begin
          ways_2_metas_97_vld <= 1'b0;
        end
        if(_zz_745) begin
          ways_2_metas_98_vld <= 1'b0;
        end
        if(_zz_746) begin
          ways_2_metas_99_vld <= 1'b0;
        end
        if(_zz_747) begin
          ways_2_metas_100_vld <= 1'b0;
        end
        if(_zz_748) begin
          ways_2_metas_101_vld <= 1'b0;
        end
        if(_zz_749) begin
          ways_2_metas_102_vld <= 1'b0;
        end
        if(_zz_750) begin
          ways_2_metas_103_vld <= 1'b0;
        end
        if(_zz_751) begin
          ways_2_metas_104_vld <= 1'b0;
        end
        if(_zz_752) begin
          ways_2_metas_105_vld <= 1'b0;
        end
        if(_zz_753) begin
          ways_2_metas_106_vld <= 1'b0;
        end
        if(_zz_754) begin
          ways_2_metas_107_vld <= 1'b0;
        end
        if(_zz_755) begin
          ways_2_metas_108_vld <= 1'b0;
        end
        if(_zz_756) begin
          ways_2_metas_109_vld <= 1'b0;
        end
        if(_zz_757) begin
          ways_2_metas_110_vld <= 1'b0;
        end
        if(_zz_758) begin
          ways_2_metas_111_vld <= 1'b0;
        end
        if(_zz_759) begin
          ways_2_metas_112_vld <= 1'b0;
        end
        if(_zz_760) begin
          ways_2_metas_113_vld <= 1'b0;
        end
        if(_zz_761) begin
          ways_2_metas_114_vld <= 1'b0;
        end
        if(_zz_762) begin
          ways_2_metas_115_vld <= 1'b0;
        end
        if(_zz_763) begin
          ways_2_metas_116_vld <= 1'b0;
        end
        if(_zz_764) begin
          ways_2_metas_117_vld <= 1'b0;
        end
        if(_zz_765) begin
          ways_2_metas_118_vld <= 1'b0;
        end
        if(_zz_766) begin
          ways_2_metas_119_vld <= 1'b0;
        end
        if(_zz_767) begin
          ways_2_metas_120_vld <= 1'b0;
        end
        if(_zz_768) begin
          ways_2_metas_121_vld <= 1'b0;
        end
        if(_zz_769) begin
          ways_2_metas_122_vld <= 1'b0;
        end
        if(_zz_770) begin
          ways_2_metas_123_vld <= 1'b0;
        end
        if(_zz_771) begin
          ways_2_metas_124_vld <= 1'b0;
        end
        if(_zz_772) begin
          ways_2_metas_125_vld <= 1'b0;
        end
        if(_zz_773) begin
          ways_2_metas_126_vld <= 1'b0;
        end
        if(_zz_774) begin
          ways_2_metas_127_vld <= 1'b0;
        end
      end else begin
        if(when_DCache_l217_2) begin
          if(cache_hit_2) begin
            if(_zz_518) begin
              ways_2_metas_0_mru <= 1'b1;
            end
            if(_zz_519) begin
              ways_2_metas_1_mru <= 1'b1;
            end
            if(_zz_520) begin
              ways_2_metas_2_mru <= 1'b1;
            end
            if(_zz_521) begin
              ways_2_metas_3_mru <= 1'b1;
            end
            if(_zz_522) begin
              ways_2_metas_4_mru <= 1'b1;
            end
            if(_zz_523) begin
              ways_2_metas_5_mru <= 1'b1;
            end
            if(_zz_524) begin
              ways_2_metas_6_mru <= 1'b1;
            end
            if(_zz_525) begin
              ways_2_metas_7_mru <= 1'b1;
            end
            if(_zz_526) begin
              ways_2_metas_8_mru <= 1'b1;
            end
            if(_zz_527) begin
              ways_2_metas_9_mru <= 1'b1;
            end
            if(_zz_528) begin
              ways_2_metas_10_mru <= 1'b1;
            end
            if(_zz_529) begin
              ways_2_metas_11_mru <= 1'b1;
            end
            if(_zz_530) begin
              ways_2_metas_12_mru <= 1'b1;
            end
            if(_zz_531) begin
              ways_2_metas_13_mru <= 1'b1;
            end
            if(_zz_532) begin
              ways_2_metas_14_mru <= 1'b1;
            end
            if(_zz_533) begin
              ways_2_metas_15_mru <= 1'b1;
            end
            if(_zz_534) begin
              ways_2_metas_16_mru <= 1'b1;
            end
            if(_zz_535) begin
              ways_2_metas_17_mru <= 1'b1;
            end
            if(_zz_536) begin
              ways_2_metas_18_mru <= 1'b1;
            end
            if(_zz_537) begin
              ways_2_metas_19_mru <= 1'b1;
            end
            if(_zz_538) begin
              ways_2_metas_20_mru <= 1'b1;
            end
            if(_zz_539) begin
              ways_2_metas_21_mru <= 1'b1;
            end
            if(_zz_540) begin
              ways_2_metas_22_mru <= 1'b1;
            end
            if(_zz_541) begin
              ways_2_metas_23_mru <= 1'b1;
            end
            if(_zz_542) begin
              ways_2_metas_24_mru <= 1'b1;
            end
            if(_zz_543) begin
              ways_2_metas_25_mru <= 1'b1;
            end
            if(_zz_544) begin
              ways_2_metas_26_mru <= 1'b1;
            end
            if(_zz_545) begin
              ways_2_metas_27_mru <= 1'b1;
            end
            if(_zz_546) begin
              ways_2_metas_28_mru <= 1'b1;
            end
            if(_zz_547) begin
              ways_2_metas_29_mru <= 1'b1;
            end
            if(_zz_548) begin
              ways_2_metas_30_mru <= 1'b1;
            end
            if(_zz_549) begin
              ways_2_metas_31_mru <= 1'b1;
            end
            if(_zz_550) begin
              ways_2_metas_32_mru <= 1'b1;
            end
            if(_zz_551) begin
              ways_2_metas_33_mru <= 1'b1;
            end
            if(_zz_552) begin
              ways_2_metas_34_mru <= 1'b1;
            end
            if(_zz_553) begin
              ways_2_metas_35_mru <= 1'b1;
            end
            if(_zz_554) begin
              ways_2_metas_36_mru <= 1'b1;
            end
            if(_zz_555) begin
              ways_2_metas_37_mru <= 1'b1;
            end
            if(_zz_556) begin
              ways_2_metas_38_mru <= 1'b1;
            end
            if(_zz_557) begin
              ways_2_metas_39_mru <= 1'b1;
            end
            if(_zz_558) begin
              ways_2_metas_40_mru <= 1'b1;
            end
            if(_zz_559) begin
              ways_2_metas_41_mru <= 1'b1;
            end
            if(_zz_560) begin
              ways_2_metas_42_mru <= 1'b1;
            end
            if(_zz_561) begin
              ways_2_metas_43_mru <= 1'b1;
            end
            if(_zz_562) begin
              ways_2_metas_44_mru <= 1'b1;
            end
            if(_zz_563) begin
              ways_2_metas_45_mru <= 1'b1;
            end
            if(_zz_564) begin
              ways_2_metas_46_mru <= 1'b1;
            end
            if(_zz_565) begin
              ways_2_metas_47_mru <= 1'b1;
            end
            if(_zz_566) begin
              ways_2_metas_48_mru <= 1'b1;
            end
            if(_zz_567) begin
              ways_2_metas_49_mru <= 1'b1;
            end
            if(_zz_568) begin
              ways_2_metas_50_mru <= 1'b1;
            end
            if(_zz_569) begin
              ways_2_metas_51_mru <= 1'b1;
            end
            if(_zz_570) begin
              ways_2_metas_52_mru <= 1'b1;
            end
            if(_zz_571) begin
              ways_2_metas_53_mru <= 1'b1;
            end
            if(_zz_572) begin
              ways_2_metas_54_mru <= 1'b1;
            end
            if(_zz_573) begin
              ways_2_metas_55_mru <= 1'b1;
            end
            if(_zz_574) begin
              ways_2_metas_56_mru <= 1'b1;
            end
            if(_zz_575) begin
              ways_2_metas_57_mru <= 1'b1;
            end
            if(_zz_576) begin
              ways_2_metas_58_mru <= 1'b1;
            end
            if(_zz_577) begin
              ways_2_metas_59_mru <= 1'b1;
            end
            if(_zz_578) begin
              ways_2_metas_60_mru <= 1'b1;
            end
            if(_zz_579) begin
              ways_2_metas_61_mru <= 1'b1;
            end
            if(_zz_580) begin
              ways_2_metas_62_mru <= 1'b1;
            end
            if(_zz_581) begin
              ways_2_metas_63_mru <= 1'b1;
            end
            if(_zz_582) begin
              ways_2_metas_64_mru <= 1'b1;
            end
            if(_zz_583) begin
              ways_2_metas_65_mru <= 1'b1;
            end
            if(_zz_584) begin
              ways_2_metas_66_mru <= 1'b1;
            end
            if(_zz_585) begin
              ways_2_metas_67_mru <= 1'b1;
            end
            if(_zz_586) begin
              ways_2_metas_68_mru <= 1'b1;
            end
            if(_zz_587) begin
              ways_2_metas_69_mru <= 1'b1;
            end
            if(_zz_588) begin
              ways_2_metas_70_mru <= 1'b1;
            end
            if(_zz_589) begin
              ways_2_metas_71_mru <= 1'b1;
            end
            if(_zz_590) begin
              ways_2_metas_72_mru <= 1'b1;
            end
            if(_zz_591) begin
              ways_2_metas_73_mru <= 1'b1;
            end
            if(_zz_592) begin
              ways_2_metas_74_mru <= 1'b1;
            end
            if(_zz_593) begin
              ways_2_metas_75_mru <= 1'b1;
            end
            if(_zz_594) begin
              ways_2_metas_76_mru <= 1'b1;
            end
            if(_zz_595) begin
              ways_2_metas_77_mru <= 1'b1;
            end
            if(_zz_596) begin
              ways_2_metas_78_mru <= 1'b1;
            end
            if(_zz_597) begin
              ways_2_metas_79_mru <= 1'b1;
            end
            if(_zz_598) begin
              ways_2_metas_80_mru <= 1'b1;
            end
            if(_zz_599) begin
              ways_2_metas_81_mru <= 1'b1;
            end
            if(_zz_600) begin
              ways_2_metas_82_mru <= 1'b1;
            end
            if(_zz_601) begin
              ways_2_metas_83_mru <= 1'b1;
            end
            if(_zz_602) begin
              ways_2_metas_84_mru <= 1'b1;
            end
            if(_zz_603) begin
              ways_2_metas_85_mru <= 1'b1;
            end
            if(_zz_604) begin
              ways_2_metas_86_mru <= 1'b1;
            end
            if(_zz_605) begin
              ways_2_metas_87_mru <= 1'b1;
            end
            if(_zz_606) begin
              ways_2_metas_88_mru <= 1'b1;
            end
            if(_zz_607) begin
              ways_2_metas_89_mru <= 1'b1;
            end
            if(_zz_608) begin
              ways_2_metas_90_mru <= 1'b1;
            end
            if(_zz_609) begin
              ways_2_metas_91_mru <= 1'b1;
            end
            if(_zz_610) begin
              ways_2_metas_92_mru <= 1'b1;
            end
            if(_zz_611) begin
              ways_2_metas_93_mru <= 1'b1;
            end
            if(_zz_612) begin
              ways_2_metas_94_mru <= 1'b1;
            end
            if(_zz_613) begin
              ways_2_metas_95_mru <= 1'b1;
            end
            if(_zz_614) begin
              ways_2_metas_96_mru <= 1'b1;
            end
            if(_zz_615) begin
              ways_2_metas_97_mru <= 1'b1;
            end
            if(_zz_616) begin
              ways_2_metas_98_mru <= 1'b1;
            end
            if(_zz_617) begin
              ways_2_metas_99_mru <= 1'b1;
            end
            if(_zz_618) begin
              ways_2_metas_100_mru <= 1'b1;
            end
            if(_zz_619) begin
              ways_2_metas_101_mru <= 1'b1;
            end
            if(_zz_620) begin
              ways_2_metas_102_mru <= 1'b1;
            end
            if(_zz_621) begin
              ways_2_metas_103_mru <= 1'b1;
            end
            if(_zz_622) begin
              ways_2_metas_104_mru <= 1'b1;
            end
            if(_zz_623) begin
              ways_2_metas_105_mru <= 1'b1;
            end
            if(_zz_624) begin
              ways_2_metas_106_mru <= 1'b1;
            end
            if(_zz_625) begin
              ways_2_metas_107_mru <= 1'b1;
            end
            if(_zz_626) begin
              ways_2_metas_108_mru <= 1'b1;
            end
            if(_zz_627) begin
              ways_2_metas_109_mru <= 1'b1;
            end
            if(_zz_628) begin
              ways_2_metas_110_mru <= 1'b1;
            end
            if(_zz_629) begin
              ways_2_metas_111_mru <= 1'b1;
            end
            if(_zz_630) begin
              ways_2_metas_112_mru <= 1'b1;
            end
            if(_zz_631) begin
              ways_2_metas_113_mru <= 1'b1;
            end
            if(_zz_632) begin
              ways_2_metas_114_mru <= 1'b1;
            end
            if(_zz_633) begin
              ways_2_metas_115_mru <= 1'b1;
            end
            if(_zz_634) begin
              ways_2_metas_116_mru <= 1'b1;
            end
            if(_zz_635) begin
              ways_2_metas_117_mru <= 1'b1;
            end
            if(_zz_636) begin
              ways_2_metas_118_mru <= 1'b1;
            end
            if(_zz_637) begin
              ways_2_metas_119_mru <= 1'b1;
            end
            if(_zz_638) begin
              ways_2_metas_120_mru <= 1'b1;
            end
            if(_zz_639) begin
              ways_2_metas_121_mru <= 1'b1;
            end
            if(_zz_640) begin
              ways_2_metas_122_mru <= 1'b1;
            end
            if(_zz_641) begin
              ways_2_metas_123_mru <= 1'b1;
            end
            if(_zz_642) begin
              ways_2_metas_124_mru <= 1'b1;
            end
            if(_zz_643) begin
              ways_2_metas_125_mru <= 1'b1;
            end
            if(_zz_644) begin
              ways_2_metas_126_mru <= 1'b1;
            end
            if(_zz_645) begin
              ways_2_metas_127_mru <= 1'b1;
            end
          end else begin
            if(_zz_518) begin
              ways_2_metas_0_mru <= 1'b0;
            end
            if(_zz_519) begin
              ways_2_metas_1_mru <= 1'b0;
            end
            if(_zz_520) begin
              ways_2_metas_2_mru <= 1'b0;
            end
            if(_zz_521) begin
              ways_2_metas_3_mru <= 1'b0;
            end
            if(_zz_522) begin
              ways_2_metas_4_mru <= 1'b0;
            end
            if(_zz_523) begin
              ways_2_metas_5_mru <= 1'b0;
            end
            if(_zz_524) begin
              ways_2_metas_6_mru <= 1'b0;
            end
            if(_zz_525) begin
              ways_2_metas_7_mru <= 1'b0;
            end
            if(_zz_526) begin
              ways_2_metas_8_mru <= 1'b0;
            end
            if(_zz_527) begin
              ways_2_metas_9_mru <= 1'b0;
            end
            if(_zz_528) begin
              ways_2_metas_10_mru <= 1'b0;
            end
            if(_zz_529) begin
              ways_2_metas_11_mru <= 1'b0;
            end
            if(_zz_530) begin
              ways_2_metas_12_mru <= 1'b0;
            end
            if(_zz_531) begin
              ways_2_metas_13_mru <= 1'b0;
            end
            if(_zz_532) begin
              ways_2_metas_14_mru <= 1'b0;
            end
            if(_zz_533) begin
              ways_2_metas_15_mru <= 1'b0;
            end
            if(_zz_534) begin
              ways_2_metas_16_mru <= 1'b0;
            end
            if(_zz_535) begin
              ways_2_metas_17_mru <= 1'b0;
            end
            if(_zz_536) begin
              ways_2_metas_18_mru <= 1'b0;
            end
            if(_zz_537) begin
              ways_2_metas_19_mru <= 1'b0;
            end
            if(_zz_538) begin
              ways_2_metas_20_mru <= 1'b0;
            end
            if(_zz_539) begin
              ways_2_metas_21_mru <= 1'b0;
            end
            if(_zz_540) begin
              ways_2_metas_22_mru <= 1'b0;
            end
            if(_zz_541) begin
              ways_2_metas_23_mru <= 1'b0;
            end
            if(_zz_542) begin
              ways_2_metas_24_mru <= 1'b0;
            end
            if(_zz_543) begin
              ways_2_metas_25_mru <= 1'b0;
            end
            if(_zz_544) begin
              ways_2_metas_26_mru <= 1'b0;
            end
            if(_zz_545) begin
              ways_2_metas_27_mru <= 1'b0;
            end
            if(_zz_546) begin
              ways_2_metas_28_mru <= 1'b0;
            end
            if(_zz_547) begin
              ways_2_metas_29_mru <= 1'b0;
            end
            if(_zz_548) begin
              ways_2_metas_30_mru <= 1'b0;
            end
            if(_zz_549) begin
              ways_2_metas_31_mru <= 1'b0;
            end
            if(_zz_550) begin
              ways_2_metas_32_mru <= 1'b0;
            end
            if(_zz_551) begin
              ways_2_metas_33_mru <= 1'b0;
            end
            if(_zz_552) begin
              ways_2_metas_34_mru <= 1'b0;
            end
            if(_zz_553) begin
              ways_2_metas_35_mru <= 1'b0;
            end
            if(_zz_554) begin
              ways_2_metas_36_mru <= 1'b0;
            end
            if(_zz_555) begin
              ways_2_metas_37_mru <= 1'b0;
            end
            if(_zz_556) begin
              ways_2_metas_38_mru <= 1'b0;
            end
            if(_zz_557) begin
              ways_2_metas_39_mru <= 1'b0;
            end
            if(_zz_558) begin
              ways_2_metas_40_mru <= 1'b0;
            end
            if(_zz_559) begin
              ways_2_metas_41_mru <= 1'b0;
            end
            if(_zz_560) begin
              ways_2_metas_42_mru <= 1'b0;
            end
            if(_zz_561) begin
              ways_2_metas_43_mru <= 1'b0;
            end
            if(_zz_562) begin
              ways_2_metas_44_mru <= 1'b0;
            end
            if(_zz_563) begin
              ways_2_metas_45_mru <= 1'b0;
            end
            if(_zz_564) begin
              ways_2_metas_46_mru <= 1'b0;
            end
            if(_zz_565) begin
              ways_2_metas_47_mru <= 1'b0;
            end
            if(_zz_566) begin
              ways_2_metas_48_mru <= 1'b0;
            end
            if(_zz_567) begin
              ways_2_metas_49_mru <= 1'b0;
            end
            if(_zz_568) begin
              ways_2_metas_50_mru <= 1'b0;
            end
            if(_zz_569) begin
              ways_2_metas_51_mru <= 1'b0;
            end
            if(_zz_570) begin
              ways_2_metas_52_mru <= 1'b0;
            end
            if(_zz_571) begin
              ways_2_metas_53_mru <= 1'b0;
            end
            if(_zz_572) begin
              ways_2_metas_54_mru <= 1'b0;
            end
            if(_zz_573) begin
              ways_2_metas_55_mru <= 1'b0;
            end
            if(_zz_574) begin
              ways_2_metas_56_mru <= 1'b0;
            end
            if(_zz_575) begin
              ways_2_metas_57_mru <= 1'b0;
            end
            if(_zz_576) begin
              ways_2_metas_58_mru <= 1'b0;
            end
            if(_zz_577) begin
              ways_2_metas_59_mru <= 1'b0;
            end
            if(_zz_578) begin
              ways_2_metas_60_mru <= 1'b0;
            end
            if(_zz_579) begin
              ways_2_metas_61_mru <= 1'b0;
            end
            if(_zz_580) begin
              ways_2_metas_62_mru <= 1'b0;
            end
            if(_zz_581) begin
              ways_2_metas_63_mru <= 1'b0;
            end
            if(_zz_582) begin
              ways_2_metas_64_mru <= 1'b0;
            end
            if(_zz_583) begin
              ways_2_metas_65_mru <= 1'b0;
            end
            if(_zz_584) begin
              ways_2_metas_66_mru <= 1'b0;
            end
            if(_zz_585) begin
              ways_2_metas_67_mru <= 1'b0;
            end
            if(_zz_586) begin
              ways_2_metas_68_mru <= 1'b0;
            end
            if(_zz_587) begin
              ways_2_metas_69_mru <= 1'b0;
            end
            if(_zz_588) begin
              ways_2_metas_70_mru <= 1'b0;
            end
            if(_zz_589) begin
              ways_2_metas_71_mru <= 1'b0;
            end
            if(_zz_590) begin
              ways_2_metas_72_mru <= 1'b0;
            end
            if(_zz_591) begin
              ways_2_metas_73_mru <= 1'b0;
            end
            if(_zz_592) begin
              ways_2_metas_74_mru <= 1'b0;
            end
            if(_zz_593) begin
              ways_2_metas_75_mru <= 1'b0;
            end
            if(_zz_594) begin
              ways_2_metas_76_mru <= 1'b0;
            end
            if(_zz_595) begin
              ways_2_metas_77_mru <= 1'b0;
            end
            if(_zz_596) begin
              ways_2_metas_78_mru <= 1'b0;
            end
            if(_zz_597) begin
              ways_2_metas_79_mru <= 1'b0;
            end
            if(_zz_598) begin
              ways_2_metas_80_mru <= 1'b0;
            end
            if(_zz_599) begin
              ways_2_metas_81_mru <= 1'b0;
            end
            if(_zz_600) begin
              ways_2_metas_82_mru <= 1'b0;
            end
            if(_zz_601) begin
              ways_2_metas_83_mru <= 1'b0;
            end
            if(_zz_602) begin
              ways_2_metas_84_mru <= 1'b0;
            end
            if(_zz_603) begin
              ways_2_metas_85_mru <= 1'b0;
            end
            if(_zz_604) begin
              ways_2_metas_86_mru <= 1'b0;
            end
            if(_zz_605) begin
              ways_2_metas_87_mru <= 1'b0;
            end
            if(_zz_606) begin
              ways_2_metas_88_mru <= 1'b0;
            end
            if(_zz_607) begin
              ways_2_metas_89_mru <= 1'b0;
            end
            if(_zz_608) begin
              ways_2_metas_90_mru <= 1'b0;
            end
            if(_zz_609) begin
              ways_2_metas_91_mru <= 1'b0;
            end
            if(_zz_610) begin
              ways_2_metas_92_mru <= 1'b0;
            end
            if(_zz_611) begin
              ways_2_metas_93_mru <= 1'b0;
            end
            if(_zz_612) begin
              ways_2_metas_94_mru <= 1'b0;
            end
            if(_zz_613) begin
              ways_2_metas_95_mru <= 1'b0;
            end
            if(_zz_614) begin
              ways_2_metas_96_mru <= 1'b0;
            end
            if(_zz_615) begin
              ways_2_metas_97_mru <= 1'b0;
            end
            if(_zz_616) begin
              ways_2_metas_98_mru <= 1'b0;
            end
            if(_zz_617) begin
              ways_2_metas_99_mru <= 1'b0;
            end
            if(_zz_618) begin
              ways_2_metas_100_mru <= 1'b0;
            end
            if(_zz_619) begin
              ways_2_metas_101_mru <= 1'b0;
            end
            if(_zz_620) begin
              ways_2_metas_102_mru <= 1'b0;
            end
            if(_zz_621) begin
              ways_2_metas_103_mru <= 1'b0;
            end
            if(_zz_622) begin
              ways_2_metas_104_mru <= 1'b0;
            end
            if(_zz_623) begin
              ways_2_metas_105_mru <= 1'b0;
            end
            if(_zz_624) begin
              ways_2_metas_106_mru <= 1'b0;
            end
            if(_zz_625) begin
              ways_2_metas_107_mru <= 1'b0;
            end
            if(_zz_626) begin
              ways_2_metas_108_mru <= 1'b0;
            end
            if(_zz_627) begin
              ways_2_metas_109_mru <= 1'b0;
            end
            if(_zz_628) begin
              ways_2_metas_110_mru <= 1'b0;
            end
            if(_zz_629) begin
              ways_2_metas_111_mru <= 1'b0;
            end
            if(_zz_630) begin
              ways_2_metas_112_mru <= 1'b0;
            end
            if(_zz_631) begin
              ways_2_metas_113_mru <= 1'b0;
            end
            if(_zz_632) begin
              ways_2_metas_114_mru <= 1'b0;
            end
            if(_zz_633) begin
              ways_2_metas_115_mru <= 1'b0;
            end
            if(_zz_634) begin
              ways_2_metas_116_mru <= 1'b0;
            end
            if(_zz_635) begin
              ways_2_metas_117_mru <= 1'b0;
            end
            if(_zz_636) begin
              ways_2_metas_118_mru <= 1'b0;
            end
            if(_zz_637) begin
              ways_2_metas_119_mru <= 1'b0;
            end
            if(_zz_638) begin
              ways_2_metas_120_mru <= 1'b0;
            end
            if(_zz_639) begin
              ways_2_metas_121_mru <= 1'b0;
            end
            if(_zz_640) begin
              ways_2_metas_122_mru <= 1'b0;
            end
            if(_zz_641) begin
              ways_2_metas_123_mru <= 1'b0;
            end
            if(_zz_642) begin
              ways_2_metas_124_mru <= 1'b0;
            end
            if(_zz_643) begin
              ways_2_metas_125_mru <= 1'b0;
            end
            if(_zz_644) begin
              ways_2_metas_126_mru <= 1'b0;
            end
            if(_zz_645) begin
              ways_2_metas_127_mru <= 1'b0;
            end
          end
        end else begin
          if(when_DCache_l224_2) begin
            if(_zz_518) begin
              ways_2_metas_0_mru <= 1'b1;
            end
            if(_zz_519) begin
              ways_2_metas_1_mru <= 1'b1;
            end
            if(_zz_520) begin
              ways_2_metas_2_mru <= 1'b1;
            end
            if(_zz_521) begin
              ways_2_metas_3_mru <= 1'b1;
            end
            if(_zz_522) begin
              ways_2_metas_4_mru <= 1'b1;
            end
            if(_zz_523) begin
              ways_2_metas_5_mru <= 1'b1;
            end
            if(_zz_524) begin
              ways_2_metas_6_mru <= 1'b1;
            end
            if(_zz_525) begin
              ways_2_metas_7_mru <= 1'b1;
            end
            if(_zz_526) begin
              ways_2_metas_8_mru <= 1'b1;
            end
            if(_zz_527) begin
              ways_2_metas_9_mru <= 1'b1;
            end
            if(_zz_528) begin
              ways_2_metas_10_mru <= 1'b1;
            end
            if(_zz_529) begin
              ways_2_metas_11_mru <= 1'b1;
            end
            if(_zz_530) begin
              ways_2_metas_12_mru <= 1'b1;
            end
            if(_zz_531) begin
              ways_2_metas_13_mru <= 1'b1;
            end
            if(_zz_532) begin
              ways_2_metas_14_mru <= 1'b1;
            end
            if(_zz_533) begin
              ways_2_metas_15_mru <= 1'b1;
            end
            if(_zz_534) begin
              ways_2_metas_16_mru <= 1'b1;
            end
            if(_zz_535) begin
              ways_2_metas_17_mru <= 1'b1;
            end
            if(_zz_536) begin
              ways_2_metas_18_mru <= 1'b1;
            end
            if(_zz_537) begin
              ways_2_metas_19_mru <= 1'b1;
            end
            if(_zz_538) begin
              ways_2_metas_20_mru <= 1'b1;
            end
            if(_zz_539) begin
              ways_2_metas_21_mru <= 1'b1;
            end
            if(_zz_540) begin
              ways_2_metas_22_mru <= 1'b1;
            end
            if(_zz_541) begin
              ways_2_metas_23_mru <= 1'b1;
            end
            if(_zz_542) begin
              ways_2_metas_24_mru <= 1'b1;
            end
            if(_zz_543) begin
              ways_2_metas_25_mru <= 1'b1;
            end
            if(_zz_544) begin
              ways_2_metas_26_mru <= 1'b1;
            end
            if(_zz_545) begin
              ways_2_metas_27_mru <= 1'b1;
            end
            if(_zz_546) begin
              ways_2_metas_28_mru <= 1'b1;
            end
            if(_zz_547) begin
              ways_2_metas_29_mru <= 1'b1;
            end
            if(_zz_548) begin
              ways_2_metas_30_mru <= 1'b1;
            end
            if(_zz_549) begin
              ways_2_metas_31_mru <= 1'b1;
            end
            if(_zz_550) begin
              ways_2_metas_32_mru <= 1'b1;
            end
            if(_zz_551) begin
              ways_2_metas_33_mru <= 1'b1;
            end
            if(_zz_552) begin
              ways_2_metas_34_mru <= 1'b1;
            end
            if(_zz_553) begin
              ways_2_metas_35_mru <= 1'b1;
            end
            if(_zz_554) begin
              ways_2_metas_36_mru <= 1'b1;
            end
            if(_zz_555) begin
              ways_2_metas_37_mru <= 1'b1;
            end
            if(_zz_556) begin
              ways_2_metas_38_mru <= 1'b1;
            end
            if(_zz_557) begin
              ways_2_metas_39_mru <= 1'b1;
            end
            if(_zz_558) begin
              ways_2_metas_40_mru <= 1'b1;
            end
            if(_zz_559) begin
              ways_2_metas_41_mru <= 1'b1;
            end
            if(_zz_560) begin
              ways_2_metas_42_mru <= 1'b1;
            end
            if(_zz_561) begin
              ways_2_metas_43_mru <= 1'b1;
            end
            if(_zz_562) begin
              ways_2_metas_44_mru <= 1'b1;
            end
            if(_zz_563) begin
              ways_2_metas_45_mru <= 1'b1;
            end
            if(_zz_564) begin
              ways_2_metas_46_mru <= 1'b1;
            end
            if(_zz_565) begin
              ways_2_metas_47_mru <= 1'b1;
            end
            if(_zz_566) begin
              ways_2_metas_48_mru <= 1'b1;
            end
            if(_zz_567) begin
              ways_2_metas_49_mru <= 1'b1;
            end
            if(_zz_568) begin
              ways_2_metas_50_mru <= 1'b1;
            end
            if(_zz_569) begin
              ways_2_metas_51_mru <= 1'b1;
            end
            if(_zz_570) begin
              ways_2_metas_52_mru <= 1'b1;
            end
            if(_zz_571) begin
              ways_2_metas_53_mru <= 1'b1;
            end
            if(_zz_572) begin
              ways_2_metas_54_mru <= 1'b1;
            end
            if(_zz_573) begin
              ways_2_metas_55_mru <= 1'b1;
            end
            if(_zz_574) begin
              ways_2_metas_56_mru <= 1'b1;
            end
            if(_zz_575) begin
              ways_2_metas_57_mru <= 1'b1;
            end
            if(_zz_576) begin
              ways_2_metas_58_mru <= 1'b1;
            end
            if(_zz_577) begin
              ways_2_metas_59_mru <= 1'b1;
            end
            if(_zz_578) begin
              ways_2_metas_60_mru <= 1'b1;
            end
            if(_zz_579) begin
              ways_2_metas_61_mru <= 1'b1;
            end
            if(_zz_580) begin
              ways_2_metas_62_mru <= 1'b1;
            end
            if(_zz_581) begin
              ways_2_metas_63_mru <= 1'b1;
            end
            if(_zz_582) begin
              ways_2_metas_64_mru <= 1'b1;
            end
            if(_zz_583) begin
              ways_2_metas_65_mru <= 1'b1;
            end
            if(_zz_584) begin
              ways_2_metas_66_mru <= 1'b1;
            end
            if(_zz_585) begin
              ways_2_metas_67_mru <= 1'b1;
            end
            if(_zz_586) begin
              ways_2_metas_68_mru <= 1'b1;
            end
            if(_zz_587) begin
              ways_2_metas_69_mru <= 1'b1;
            end
            if(_zz_588) begin
              ways_2_metas_70_mru <= 1'b1;
            end
            if(_zz_589) begin
              ways_2_metas_71_mru <= 1'b1;
            end
            if(_zz_590) begin
              ways_2_metas_72_mru <= 1'b1;
            end
            if(_zz_591) begin
              ways_2_metas_73_mru <= 1'b1;
            end
            if(_zz_592) begin
              ways_2_metas_74_mru <= 1'b1;
            end
            if(_zz_593) begin
              ways_2_metas_75_mru <= 1'b1;
            end
            if(_zz_594) begin
              ways_2_metas_76_mru <= 1'b1;
            end
            if(_zz_595) begin
              ways_2_metas_77_mru <= 1'b1;
            end
            if(_zz_596) begin
              ways_2_metas_78_mru <= 1'b1;
            end
            if(_zz_597) begin
              ways_2_metas_79_mru <= 1'b1;
            end
            if(_zz_598) begin
              ways_2_metas_80_mru <= 1'b1;
            end
            if(_zz_599) begin
              ways_2_metas_81_mru <= 1'b1;
            end
            if(_zz_600) begin
              ways_2_metas_82_mru <= 1'b1;
            end
            if(_zz_601) begin
              ways_2_metas_83_mru <= 1'b1;
            end
            if(_zz_602) begin
              ways_2_metas_84_mru <= 1'b1;
            end
            if(_zz_603) begin
              ways_2_metas_85_mru <= 1'b1;
            end
            if(_zz_604) begin
              ways_2_metas_86_mru <= 1'b1;
            end
            if(_zz_605) begin
              ways_2_metas_87_mru <= 1'b1;
            end
            if(_zz_606) begin
              ways_2_metas_88_mru <= 1'b1;
            end
            if(_zz_607) begin
              ways_2_metas_89_mru <= 1'b1;
            end
            if(_zz_608) begin
              ways_2_metas_90_mru <= 1'b1;
            end
            if(_zz_609) begin
              ways_2_metas_91_mru <= 1'b1;
            end
            if(_zz_610) begin
              ways_2_metas_92_mru <= 1'b1;
            end
            if(_zz_611) begin
              ways_2_metas_93_mru <= 1'b1;
            end
            if(_zz_612) begin
              ways_2_metas_94_mru <= 1'b1;
            end
            if(_zz_613) begin
              ways_2_metas_95_mru <= 1'b1;
            end
            if(_zz_614) begin
              ways_2_metas_96_mru <= 1'b1;
            end
            if(_zz_615) begin
              ways_2_metas_97_mru <= 1'b1;
            end
            if(_zz_616) begin
              ways_2_metas_98_mru <= 1'b1;
            end
            if(_zz_617) begin
              ways_2_metas_99_mru <= 1'b1;
            end
            if(_zz_618) begin
              ways_2_metas_100_mru <= 1'b1;
            end
            if(_zz_619) begin
              ways_2_metas_101_mru <= 1'b1;
            end
            if(_zz_620) begin
              ways_2_metas_102_mru <= 1'b1;
            end
            if(_zz_621) begin
              ways_2_metas_103_mru <= 1'b1;
            end
            if(_zz_622) begin
              ways_2_metas_104_mru <= 1'b1;
            end
            if(_zz_623) begin
              ways_2_metas_105_mru <= 1'b1;
            end
            if(_zz_624) begin
              ways_2_metas_106_mru <= 1'b1;
            end
            if(_zz_625) begin
              ways_2_metas_107_mru <= 1'b1;
            end
            if(_zz_626) begin
              ways_2_metas_108_mru <= 1'b1;
            end
            if(_zz_627) begin
              ways_2_metas_109_mru <= 1'b1;
            end
            if(_zz_628) begin
              ways_2_metas_110_mru <= 1'b1;
            end
            if(_zz_629) begin
              ways_2_metas_111_mru <= 1'b1;
            end
            if(_zz_630) begin
              ways_2_metas_112_mru <= 1'b1;
            end
            if(_zz_631) begin
              ways_2_metas_113_mru <= 1'b1;
            end
            if(_zz_632) begin
              ways_2_metas_114_mru <= 1'b1;
            end
            if(_zz_633) begin
              ways_2_metas_115_mru <= 1'b1;
            end
            if(_zz_634) begin
              ways_2_metas_116_mru <= 1'b1;
            end
            if(_zz_635) begin
              ways_2_metas_117_mru <= 1'b1;
            end
            if(_zz_636) begin
              ways_2_metas_118_mru <= 1'b1;
            end
            if(_zz_637) begin
              ways_2_metas_119_mru <= 1'b1;
            end
            if(_zz_638) begin
              ways_2_metas_120_mru <= 1'b1;
            end
            if(_zz_639) begin
              ways_2_metas_121_mru <= 1'b1;
            end
            if(_zz_640) begin
              ways_2_metas_122_mru <= 1'b1;
            end
            if(_zz_641) begin
              ways_2_metas_123_mru <= 1'b1;
            end
            if(_zz_642) begin
              ways_2_metas_124_mru <= 1'b1;
            end
            if(_zz_643) begin
              ways_2_metas_125_mru <= 1'b1;
            end
            if(_zz_644) begin
              ways_2_metas_126_mru <= 1'b1;
            end
            if(_zz_645) begin
              ways_2_metas_127_mru <= 1'b1;
            end
          end else begin
            if(when_DCache_l227_2) begin
              if(_zz_518) begin
                ways_2_metas_0_vld <= 1'b1;
              end
              if(_zz_519) begin
                ways_2_metas_1_vld <= 1'b1;
              end
              if(_zz_520) begin
                ways_2_metas_2_vld <= 1'b1;
              end
              if(_zz_521) begin
                ways_2_metas_3_vld <= 1'b1;
              end
              if(_zz_522) begin
                ways_2_metas_4_vld <= 1'b1;
              end
              if(_zz_523) begin
                ways_2_metas_5_vld <= 1'b1;
              end
              if(_zz_524) begin
                ways_2_metas_6_vld <= 1'b1;
              end
              if(_zz_525) begin
                ways_2_metas_7_vld <= 1'b1;
              end
              if(_zz_526) begin
                ways_2_metas_8_vld <= 1'b1;
              end
              if(_zz_527) begin
                ways_2_metas_9_vld <= 1'b1;
              end
              if(_zz_528) begin
                ways_2_metas_10_vld <= 1'b1;
              end
              if(_zz_529) begin
                ways_2_metas_11_vld <= 1'b1;
              end
              if(_zz_530) begin
                ways_2_metas_12_vld <= 1'b1;
              end
              if(_zz_531) begin
                ways_2_metas_13_vld <= 1'b1;
              end
              if(_zz_532) begin
                ways_2_metas_14_vld <= 1'b1;
              end
              if(_zz_533) begin
                ways_2_metas_15_vld <= 1'b1;
              end
              if(_zz_534) begin
                ways_2_metas_16_vld <= 1'b1;
              end
              if(_zz_535) begin
                ways_2_metas_17_vld <= 1'b1;
              end
              if(_zz_536) begin
                ways_2_metas_18_vld <= 1'b1;
              end
              if(_zz_537) begin
                ways_2_metas_19_vld <= 1'b1;
              end
              if(_zz_538) begin
                ways_2_metas_20_vld <= 1'b1;
              end
              if(_zz_539) begin
                ways_2_metas_21_vld <= 1'b1;
              end
              if(_zz_540) begin
                ways_2_metas_22_vld <= 1'b1;
              end
              if(_zz_541) begin
                ways_2_metas_23_vld <= 1'b1;
              end
              if(_zz_542) begin
                ways_2_metas_24_vld <= 1'b1;
              end
              if(_zz_543) begin
                ways_2_metas_25_vld <= 1'b1;
              end
              if(_zz_544) begin
                ways_2_metas_26_vld <= 1'b1;
              end
              if(_zz_545) begin
                ways_2_metas_27_vld <= 1'b1;
              end
              if(_zz_546) begin
                ways_2_metas_28_vld <= 1'b1;
              end
              if(_zz_547) begin
                ways_2_metas_29_vld <= 1'b1;
              end
              if(_zz_548) begin
                ways_2_metas_30_vld <= 1'b1;
              end
              if(_zz_549) begin
                ways_2_metas_31_vld <= 1'b1;
              end
              if(_zz_550) begin
                ways_2_metas_32_vld <= 1'b1;
              end
              if(_zz_551) begin
                ways_2_metas_33_vld <= 1'b1;
              end
              if(_zz_552) begin
                ways_2_metas_34_vld <= 1'b1;
              end
              if(_zz_553) begin
                ways_2_metas_35_vld <= 1'b1;
              end
              if(_zz_554) begin
                ways_2_metas_36_vld <= 1'b1;
              end
              if(_zz_555) begin
                ways_2_metas_37_vld <= 1'b1;
              end
              if(_zz_556) begin
                ways_2_metas_38_vld <= 1'b1;
              end
              if(_zz_557) begin
                ways_2_metas_39_vld <= 1'b1;
              end
              if(_zz_558) begin
                ways_2_metas_40_vld <= 1'b1;
              end
              if(_zz_559) begin
                ways_2_metas_41_vld <= 1'b1;
              end
              if(_zz_560) begin
                ways_2_metas_42_vld <= 1'b1;
              end
              if(_zz_561) begin
                ways_2_metas_43_vld <= 1'b1;
              end
              if(_zz_562) begin
                ways_2_metas_44_vld <= 1'b1;
              end
              if(_zz_563) begin
                ways_2_metas_45_vld <= 1'b1;
              end
              if(_zz_564) begin
                ways_2_metas_46_vld <= 1'b1;
              end
              if(_zz_565) begin
                ways_2_metas_47_vld <= 1'b1;
              end
              if(_zz_566) begin
                ways_2_metas_48_vld <= 1'b1;
              end
              if(_zz_567) begin
                ways_2_metas_49_vld <= 1'b1;
              end
              if(_zz_568) begin
                ways_2_metas_50_vld <= 1'b1;
              end
              if(_zz_569) begin
                ways_2_metas_51_vld <= 1'b1;
              end
              if(_zz_570) begin
                ways_2_metas_52_vld <= 1'b1;
              end
              if(_zz_571) begin
                ways_2_metas_53_vld <= 1'b1;
              end
              if(_zz_572) begin
                ways_2_metas_54_vld <= 1'b1;
              end
              if(_zz_573) begin
                ways_2_metas_55_vld <= 1'b1;
              end
              if(_zz_574) begin
                ways_2_metas_56_vld <= 1'b1;
              end
              if(_zz_575) begin
                ways_2_metas_57_vld <= 1'b1;
              end
              if(_zz_576) begin
                ways_2_metas_58_vld <= 1'b1;
              end
              if(_zz_577) begin
                ways_2_metas_59_vld <= 1'b1;
              end
              if(_zz_578) begin
                ways_2_metas_60_vld <= 1'b1;
              end
              if(_zz_579) begin
                ways_2_metas_61_vld <= 1'b1;
              end
              if(_zz_580) begin
                ways_2_metas_62_vld <= 1'b1;
              end
              if(_zz_581) begin
                ways_2_metas_63_vld <= 1'b1;
              end
              if(_zz_582) begin
                ways_2_metas_64_vld <= 1'b1;
              end
              if(_zz_583) begin
                ways_2_metas_65_vld <= 1'b1;
              end
              if(_zz_584) begin
                ways_2_metas_66_vld <= 1'b1;
              end
              if(_zz_585) begin
                ways_2_metas_67_vld <= 1'b1;
              end
              if(_zz_586) begin
                ways_2_metas_68_vld <= 1'b1;
              end
              if(_zz_587) begin
                ways_2_metas_69_vld <= 1'b1;
              end
              if(_zz_588) begin
                ways_2_metas_70_vld <= 1'b1;
              end
              if(_zz_589) begin
                ways_2_metas_71_vld <= 1'b1;
              end
              if(_zz_590) begin
                ways_2_metas_72_vld <= 1'b1;
              end
              if(_zz_591) begin
                ways_2_metas_73_vld <= 1'b1;
              end
              if(_zz_592) begin
                ways_2_metas_74_vld <= 1'b1;
              end
              if(_zz_593) begin
                ways_2_metas_75_vld <= 1'b1;
              end
              if(_zz_594) begin
                ways_2_metas_76_vld <= 1'b1;
              end
              if(_zz_595) begin
                ways_2_metas_77_vld <= 1'b1;
              end
              if(_zz_596) begin
                ways_2_metas_78_vld <= 1'b1;
              end
              if(_zz_597) begin
                ways_2_metas_79_vld <= 1'b1;
              end
              if(_zz_598) begin
                ways_2_metas_80_vld <= 1'b1;
              end
              if(_zz_599) begin
                ways_2_metas_81_vld <= 1'b1;
              end
              if(_zz_600) begin
                ways_2_metas_82_vld <= 1'b1;
              end
              if(_zz_601) begin
                ways_2_metas_83_vld <= 1'b1;
              end
              if(_zz_602) begin
                ways_2_metas_84_vld <= 1'b1;
              end
              if(_zz_603) begin
                ways_2_metas_85_vld <= 1'b1;
              end
              if(_zz_604) begin
                ways_2_metas_86_vld <= 1'b1;
              end
              if(_zz_605) begin
                ways_2_metas_87_vld <= 1'b1;
              end
              if(_zz_606) begin
                ways_2_metas_88_vld <= 1'b1;
              end
              if(_zz_607) begin
                ways_2_metas_89_vld <= 1'b1;
              end
              if(_zz_608) begin
                ways_2_metas_90_vld <= 1'b1;
              end
              if(_zz_609) begin
                ways_2_metas_91_vld <= 1'b1;
              end
              if(_zz_610) begin
                ways_2_metas_92_vld <= 1'b1;
              end
              if(_zz_611) begin
                ways_2_metas_93_vld <= 1'b1;
              end
              if(_zz_612) begin
                ways_2_metas_94_vld <= 1'b1;
              end
              if(_zz_613) begin
                ways_2_metas_95_vld <= 1'b1;
              end
              if(_zz_614) begin
                ways_2_metas_96_vld <= 1'b1;
              end
              if(_zz_615) begin
                ways_2_metas_97_vld <= 1'b1;
              end
              if(_zz_616) begin
                ways_2_metas_98_vld <= 1'b1;
              end
              if(_zz_617) begin
                ways_2_metas_99_vld <= 1'b1;
              end
              if(_zz_618) begin
                ways_2_metas_100_vld <= 1'b1;
              end
              if(_zz_619) begin
                ways_2_metas_101_vld <= 1'b1;
              end
              if(_zz_620) begin
                ways_2_metas_102_vld <= 1'b1;
              end
              if(_zz_621) begin
                ways_2_metas_103_vld <= 1'b1;
              end
              if(_zz_622) begin
                ways_2_metas_104_vld <= 1'b1;
              end
              if(_zz_623) begin
                ways_2_metas_105_vld <= 1'b1;
              end
              if(_zz_624) begin
                ways_2_metas_106_vld <= 1'b1;
              end
              if(_zz_625) begin
                ways_2_metas_107_vld <= 1'b1;
              end
              if(_zz_626) begin
                ways_2_metas_108_vld <= 1'b1;
              end
              if(_zz_627) begin
                ways_2_metas_109_vld <= 1'b1;
              end
              if(_zz_628) begin
                ways_2_metas_110_vld <= 1'b1;
              end
              if(_zz_629) begin
                ways_2_metas_111_vld <= 1'b1;
              end
              if(_zz_630) begin
                ways_2_metas_112_vld <= 1'b1;
              end
              if(_zz_631) begin
                ways_2_metas_113_vld <= 1'b1;
              end
              if(_zz_632) begin
                ways_2_metas_114_vld <= 1'b1;
              end
              if(_zz_633) begin
                ways_2_metas_115_vld <= 1'b1;
              end
              if(_zz_634) begin
                ways_2_metas_116_vld <= 1'b1;
              end
              if(_zz_635) begin
                ways_2_metas_117_vld <= 1'b1;
              end
              if(_zz_636) begin
                ways_2_metas_118_vld <= 1'b1;
              end
              if(_zz_637) begin
                ways_2_metas_119_vld <= 1'b1;
              end
              if(_zz_638) begin
                ways_2_metas_120_vld <= 1'b1;
              end
              if(_zz_639) begin
                ways_2_metas_121_vld <= 1'b1;
              end
              if(_zz_640) begin
                ways_2_metas_122_vld <= 1'b1;
              end
              if(_zz_641) begin
                ways_2_metas_123_vld <= 1'b1;
              end
              if(_zz_642) begin
                ways_2_metas_124_vld <= 1'b1;
              end
              if(_zz_643) begin
                ways_2_metas_125_vld <= 1'b1;
              end
              if(_zz_644) begin
                ways_2_metas_126_vld <= 1'b1;
              end
              if(_zz_645) begin
                ways_2_metas_127_vld <= 1'b1;
              end
            end
          end
        end
      end
      if(when_DCache_l232_2) begin
        if(_zz_518) begin
          ways_2_metas_0_tag <= cpu_tag;
        end
        if(_zz_519) begin
          ways_2_metas_1_tag <= cpu_tag;
        end
        if(_zz_520) begin
          ways_2_metas_2_tag <= cpu_tag;
        end
        if(_zz_521) begin
          ways_2_metas_3_tag <= cpu_tag;
        end
        if(_zz_522) begin
          ways_2_metas_4_tag <= cpu_tag;
        end
        if(_zz_523) begin
          ways_2_metas_5_tag <= cpu_tag;
        end
        if(_zz_524) begin
          ways_2_metas_6_tag <= cpu_tag;
        end
        if(_zz_525) begin
          ways_2_metas_7_tag <= cpu_tag;
        end
        if(_zz_526) begin
          ways_2_metas_8_tag <= cpu_tag;
        end
        if(_zz_527) begin
          ways_2_metas_9_tag <= cpu_tag;
        end
        if(_zz_528) begin
          ways_2_metas_10_tag <= cpu_tag;
        end
        if(_zz_529) begin
          ways_2_metas_11_tag <= cpu_tag;
        end
        if(_zz_530) begin
          ways_2_metas_12_tag <= cpu_tag;
        end
        if(_zz_531) begin
          ways_2_metas_13_tag <= cpu_tag;
        end
        if(_zz_532) begin
          ways_2_metas_14_tag <= cpu_tag;
        end
        if(_zz_533) begin
          ways_2_metas_15_tag <= cpu_tag;
        end
        if(_zz_534) begin
          ways_2_metas_16_tag <= cpu_tag;
        end
        if(_zz_535) begin
          ways_2_metas_17_tag <= cpu_tag;
        end
        if(_zz_536) begin
          ways_2_metas_18_tag <= cpu_tag;
        end
        if(_zz_537) begin
          ways_2_metas_19_tag <= cpu_tag;
        end
        if(_zz_538) begin
          ways_2_metas_20_tag <= cpu_tag;
        end
        if(_zz_539) begin
          ways_2_metas_21_tag <= cpu_tag;
        end
        if(_zz_540) begin
          ways_2_metas_22_tag <= cpu_tag;
        end
        if(_zz_541) begin
          ways_2_metas_23_tag <= cpu_tag;
        end
        if(_zz_542) begin
          ways_2_metas_24_tag <= cpu_tag;
        end
        if(_zz_543) begin
          ways_2_metas_25_tag <= cpu_tag;
        end
        if(_zz_544) begin
          ways_2_metas_26_tag <= cpu_tag;
        end
        if(_zz_545) begin
          ways_2_metas_27_tag <= cpu_tag;
        end
        if(_zz_546) begin
          ways_2_metas_28_tag <= cpu_tag;
        end
        if(_zz_547) begin
          ways_2_metas_29_tag <= cpu_tag;
        end
        if(_zz_548) begin
          ways_2_metas_30_tag <= cpu_tag;
        end
        if(_zz_549) begin
          ways_2_metas_31_tag <= cpu_tag;
        end
        if(_zz_550) begin
          ways_2_metas_32_tag <= cpu_tag;
        end
        if(_zz_551) begin
          ways_2_metas_33_tag <= cpu_tag;
        end
        if(_zz_552) begin
          ways_2_metas_34_tag <= cpu_tag;
        end
        if(_zz_553) begin
          ways_2_metas_35_tag <= cpu_tag;
        end
        if(_zz_554) begin
          ways_2_metas_36_tag <= cpu_tag;
        end
        if(_zz_555) begin
          ways_2_metas_37_tag <= cpu_tag;
        end
        if(_zz_556) begin
          ways_2_metas_38_tag <= cpu_tag;
        end
        if(_zz_557) begin
          ways_2_metas_39_tag <= cpu_tag;
        end
        if(_zz_558) begin
          ways_2_metas_40_tag <= cpu_tag;
        end
        if(_zz_559) begin
          ways_2_metas_41_tag <= cpu_tag;
        end
        if(_zz_560) begin
          ways_2_metas_42_tag <= cpu_tag;
        end
        if(_zz_561) begin
          ways_2_metas_43_tag <= cpu_tag;
        end
        if(_zz_562) begin
          ways_2_metas_44_tag <= cpu_tag;
        end
        if(_zz_563) begin
          ways_2_metas_45_tag <= cpu_tag;
        end
        if(_zz_564) begin
          ways_2_metas_46_tag <= cpu_tag;
        end
        if(_zz_565) begin
          ways_2_metas_47_tag <= cpu_tag;
        end
        if(_zz_566) begin
          ways_2_metas_48_tag <= cpu_tag;
        end
        if(_zz_567) begin
          ways_2_metas_49_tag <= cpu_tag;
        end
        if(_zz_568) begin
          ways_2_metas_50_tag <= cpu_tag;
        end
        if(_zz_569) begin
          ways_2_metas_51_tag <= cpu_tag;
        end
        if(_zz_570) begin
          ways_2_metas_52_tag <= cpu_tag;
        end
        if(_zz_571) begin
          ways_2_metas_53_tag <= cpu_tag;
        end
        if(_zz_572) begin
          ways_2_metas_54_tag <= cpu_tag;
        end
        if(_zz_573) begin
          ways_2_metas_55_tag <= cpu_tag;
        end
        if(_zz_574) begin
          ways_2_metas_56_tag <= cpu_tag;
        end
        if(_zz_575) begin
          ways_2_metas_57_tag <= cpu_tag;
        end
        if(_zz_576) begin
          ways_2_metas_58_tag <= cpu_tag;
        end
        if(_zz_577) begin
          ways_2_metas_59_tag <= cpu_tag;
        end
        if(_zz_578) begin
          ways_2_metas_60_tag <= cpu_tag;
        end
        if(_zz_579) begin
          ways_2_metas_61_tag <= cpu_tag;
        end
        if(_zz_580) begin
          ways_2_metas_62_tag <= cpu_tag;
        end
        if(_zz_581) begin
          ways_2_metas_63_tag <= cpu_tag;
        end
        if(_zz_582) begin
          ways_2_metas_64_tag <= cpu_tag;
        end
        if(_zz_583) begin
          ways_2_metas_65_tag <= cpu_tag;
        end
        if(_zz_584) begin
          ways_2_metas_66_tag <= cpu_tag;
        end
        if(_zz_585) begin
          ways_2_metas_67_tag <= cpu_tag;
        end
        if(_zz_586) begin
          ways_2_metas_68_tag <= cpu_tag;
        end
        if(_zz_587) begin
          ways_2_metas_69_tag <= cpu_tag;
        end
        if(_zz_588) begin
          ways_2_metas_70_tag <= cpu_tag;
        end
        if(_zz_589) begin
          ways_2_metas_71_tag <= cpu_tag;
        end
        if(_zz_590) begin
          ways_2_metas_72_tag <= cpu_tag;
        end
        if(_zz_591) begin
          ways_2_metas_73_tag <= cpu_tag;
        end
        if(_zz_592) begin
          ways_2_metas_74_tag <= cpu_tag;
        end
        if(_zz_593) begin
          ways_2_metas_75_tag <= cpu_tag;
        end
        if(_zz_594) begin
          ways_2_metas_76_tag <= cpu_tag;
        end
        if(_zz_595) begin
          ways_2_metas_77_tag <= cpu_tag;
        end
        if(_zz_596) begin
          ways_2_metas_78_tag <= cpu_tag;
        end
        if(_zz_597) begin
          ways_2_metas_79_tag <= cpu_tag;
        end
        if(_zz_598) begin
          ways_2_metas_80_tag <= cpu_tag;
        end
        if(_zz_599) begin
          ways_2_metas_81_tag <= cpu_tag;
        end
        if(_zz_600) begin
          ways_2_metas_82_tag <= cpu_tag;
        end
        if(_zz_601) begin
          ways_2_metas_83_tag <= cpu_tag;
        end
        if(_zz_602) begin
          ways_2_metas_84_tag <= cpu_tag;
        end
        if(_zz_603) begin
          ways_2_metas_85_tag <= cpu_tag;
        end
        if(_zz_604) begin
          ways_2_metas_86_tag <= cpu_tag;
        end
        if(_zz_605) begin
          ways_2_metas_87_tag <= cpu_tag;
        end
        if(_zz_606) begin
          ways_2_metas_88_tag <= cpu_tag;
        end
        if(_zz_607) begin
          ways_2_metas_89_tag <= cpu_tag;
        end
        if(_zz_608) begin
          ways_2_metas_90_tag <= cpu_tag;
        end
        if(_zz_609) begin
          ways_2_metas_91_tag <= cpu_tag;
        end
        if(_zz_610) begin
          ways_2_metas_92_tag <= cpu_tag;
        end
        if(_zz_611) begin
          ways_2_metas_93_tag <= cpu_tag;
        end
        if(_zz_612) begin
          ways_2_metas_94_tag <= cpu_tag;
        end
        if(_zz_613) begin
          ways_2_metas_95_tag <= cpu_tag;
        end
        if(_zz_614) begin
          ways_2_metas_96_tag <= cpu_tag;
        end
        if(_zz_615) begin
          ways_2_metas_97_tag <= cpu_tag;
        end
        if(_zz_616) begin
          ways_2_metas_98_tag <= cpu_tag;
        end
        if(_zz_617) begin
          ways_2_metas_99_tag <= cpu_tag;
        end
        if(_zz_618) begin
          ways_2_metas_100_tag <= cpu_tag;
        end
        if(_zz_619) begin
          ways_2_metas_101_tag <= cpu_tag;
        end
        if(_zz_620) begin
          ways_2_metas_102_tag <= cpu_tag;
        end
        if(_zz_621) begin
          ways_2_metas_103_tag <= cpu_tag;
        end
        if(_zz_622) begin
          ways_2_metas_104_tag <= cpu_tag;
        end
        if(_zz_623) begin
          ways_2_metas_105_tag <= cpu_tag;
        end
        if(_zz_624) begin
          ways_2_metas_106_tag <= cpu_tag;
        end
        if(_zz_625) begin
          ways_2_metas_107_tag <= cpu_tag;
        end
        if(_zz_626) begin
          ways_2_metas_108_tag <= cpu_tag;
        end
        if(_zz_627) begin
          ways_2_metas_109_tag <= cpu_tag;
        end
        if(_zz_628) begin
          ways_2_metas_110_tag <= cpu_tag;
        end
        if(_zz_629) begin
          ways_2_metas_111_tag <= cpu_tag;
        end
        if(_zz_630) begin
          ways_2_metas_112_tag <= cpu_tag;
        end
        if(_zz_631) begin
          ways_2_metas_113_tag <= cpu_tag;
        end
        if(_zz_632) begin
          ways_2_metas_114_tag <= cpu_tag;
        end
        if(_zz_633) begin
          ways_2_metas_115_tag <= cpu_tag;
        end
        if(_zz_634) begin
          ways_2_metas_116_tag <= cpu_tag;
        end
        if(_zz_635) begin
          ways_2_metas_117_tag <= cpu_tag;
        end
        if(_zz_636) begin
          ways_2_metas_118_tag <= cpu_tag;
        end
        if(_zz_637) begin
          ways_2_metas_119_tag <= cpu_tag;
        end
        if(_zz_638) begin
          ways_2_metas_120_tag <= cpu_tag;
        end
        if(_zz_639) begin
          ways_2_metas_121_tag <= cpu_tag;
        end
        if(_zz_640) begin
          ways_2_metas_122_tag <= cpu_tag;
        end
        if(_zz_641) begin
          ways_2_metas_123_tag <= cpu_tag;
        end
        if(_zz_642) begin
          ways_2_metas_124_tag <= cpu_tag;
        end
        if(_zz_643) begin
          ways_2_metas_125_tag <= cpu_tag;
        end
        if(_zz_644) begin
          ways_2_metas_126_tag <= cpu_tag;
        end
        if(_zz_645) begin
          ways_2_metas_127_tag <= cpu_tag;
        end
      end
      if(when_DCache_l237_2) begin
        cpu_cmd_ready_1 <= 1'b0;
      end else begin
        if(when_DCache_l240_2) begin
          cpu_cmd_ready_1 <= 1'b1;
        end
      end
      if(flush_busy) begin
        if(_zz_905) begin
          ways_3_metas_0_mru <= 1'b0;
        end
        if(_zz_906) begin
          ways_3_metas_1_mru <= 1'b0;
        end
        if(_zz_907) begin
          ways_3_metas_2_mru <= 1'b0;
        end
        if(_zz_908) begin
          ways_3_metas_3_mru <= 1'b0;
        end
        if(_zz_909) begin
          ways_3_metas_4_mru <= 1'b0;
        end
        if(_zz_910) begin
          ways_3_metas_5_mru <= 1'b0;
        end
        if(_zz_911) begin
          ways_3_metas_6_mru <= 1'b0;
        end
        if(_zz_912) begin
          ways_3_metas_7_mru <= 1'b0;
        end
        if(_zz_913) begin
          ways_3_metas_8_mru <= 1'b0;
        end
        if(_zz_914) begin
          ways_3_metas_9_mru <= 1'b0;
        end
        if(_zz_915) begin
          ways_3_metas_10_mru <= 1'b0;
        end
        if(_zz_916) begin
          ways_3_metas_11_mru <= 1'b0;
        end
        if(_zz_917) begin
          ways_3_metas_12_mru <= 1'b0;
        end
        if(_zz_918) begin
          ways_3_metas_13_mru <= 1'b0;
        end
        if(_zz_919) begin
          ways_3_metas_14_mru <= 1'b0;
        end
        if(_zz_920) begin
          ways_3_metas_15_mru <= 1'b0;
        end
        if(_zz_921) begin
          ways_3_metas_16_mru <= 1'b0;
        end
        if(_zz_922) begin
          ways_3_metas_17_mru <= 1'b0;
        end
        if(_zz_923) begin
          ways_3_metas_18_mru <= 1'b0;
        end
        if(_zz_924) begin
          ways_3_metas_19_mru <= 1'b0;
        end
        if(_zz_925) begin
          ways_3_metas_20_mru <= 1'b0;
        end
        if(_zz_926) begin
          ways_3_metas_21_mru <= 1'b0;
        end
        if(_zz_927) begin
          ways_3_metas_22_mru <= 1'b0;
        end
        if(_zz_928) begin
          ways_3_metas_23_mru <= 1'b0;
        end
        if(_zz_929) begin
          ways_3_metas_24_mru <= 1'b0;
        end
        if(_zz_930) begin
          ways_3_metas_25_mru <= 1'b0;
        end
        if(_zz_931) begin
          ways_3_metas_26_mru <= 1'b0;
        end
        if(_zz_932) begin
          ways_3_metas_27_mru <= 1'b0;
        end
        if(_zz_933) begin
          ways_3_metas_28_mru <= 1'b0;
        end
        if(_zz_934) begin
          ways_3_metas_29_mru <= 1'b0;
        end
        if(_zz_935) begin
          ways_3_metas_30_mru <= 1'b0;
        end
        if(_zz_936) begin
          ways_3_metas_31_mru <= 1'b0;
        end
        if(_zz_937) begin
          ways_3_metas_32_mru <= 1'b0;
        end
        if(_zz_938) begin
          ways_3_metas_33_mru <= 1'b0;
        end
        if(_zz_939) begin
          ways_3_metas_34_mru <= 1'b0;
        end
        if(_zz_940) begin
          ways_3_metas_35_mru <= 1'b0;
        end
        if(_zz_941) begin
          ways_3_metas_36_mru <= 1'b0;
        end
        if(_zz_942) begin
          ways_3_metas_37_mru <= 1'b0;
        end
        if(_zz_943) begin
          ways_3_metas_38_mru <= 1'b0;
        end
        if(_zz_944) begin
          ways_3_metas_39_mru <= 1'b0;
        end
        if(_zz_945) begin
          ways_3_metas_40_mru <= 1'b0;
        end
        if(_zz_946) begin
          ways_3_metas_41_mru <= 1'b0;
        end
        if(_zz_947) begin
          ways_3_metas_42_mru <= 1'b0;
        end
        if(_zz_948) begin
          ways_3_metas_43_mru <= 1'b0;
        end
        if(_zz_949) begin
          ways_3_metas_44_mru <= 1'b0;
        end
        if(_zz_950) begin
          ways_3_metas_45_mru <= 1'b0;
        end
        if(_zz_951) begin
          ways_3_metas_46_mru <= 1'b0;
        end
        if(_zz_952) begin
          ways_3_metas_47_mru <= 1'b0;
        end
        if(_zz_953) begin
          ways_3_metas_48_mru <= 1'b0;
        end
        if(_zz_954) begin
          ways_3_metas_49_mru <= 1'b0;
        end
        if(_zz_955) begin
          ways_3_metas_50_mru <= 1'b0;
        end
        if(_zz_956) begin
          ways_3_metas_51_mru <= 1'b0;
        end
        if(_zz_957) begin
          ways_3_metas_52_mru <= 1'b0;
        end
        if(_zz_958) begin
          ways_3_metas_53_mru <= 1'b0;
        end
        if(_zz_959) begin
          ways_3_metas_54_mru <= 1'b0;
        end
        if(_zz_960) begin
          ways_3_metas_55_mru <= 1'b0;
        end
        if(_zz_961) begin
          ways_3_metas_56_mru <= 1'b0;
        end
        if(_zz_962) begin
          ways_3_metas_57_mru <= 1'b0;
        end
        if(_zz_963) begin
          ways_3_metas_58_mru <= 1'b0;
        end
        if(_zz_964) begin
          ways_3_metas_59_mru <= 1'b0;
        end
        if(_zz_965) begin
          ways_3_metas_60_mru <= 1'b0;
        end
        if(_zz_966) begin
          ways_3_metas_61_mru <= 1'b0;
        end
        if(_zz_967) begin
          ways_3_metas_62_mru <= 1'b0;
        end
        if(_zz_968) begin
          ways_3_metas_63_mru <= 1'b0;
        end
        if(_zz_969) begin
          ways_3_metas_64_mru <= 1'b0;
        end
        if(_zz_970) begin
          ways_3_metas_65_mru <= 1'b0;
        end
        if(_zz_971) begin
          ways_3_metas_66_mru <= 1'b0;
        end
        if(_zz_972) begin
          ways_3_metas_67_mru <= 1'b0;
        end
        if(_zz_973) begin
          ways_3_metas_68_mru <= 1'b0;
        end
        if(_zz_974) begin
          ways_3_metas_69_mru <= 1'b0;
        end
        if(_zz_975) begin
          ways_3_metas_70_mru <= 1'b0;
        end
        if(_zz_976) begin
          ways_3_metas_71_mru <= 1'b0;
        end
        if(_zz_977) begin
          ways_3_metas_72_mru <= 1'b0;
        end
        if(_zz_978) begin
          ways_3_metas_73_mru <= 1'b0;
        end
        if(_zz_979) begin
          ways_3_metas_74_mru <= 1'b0;
        end
        if(_zz_980) begin
          ways_3_metas_75_mru <= 1'b0;
        end
        if(_zz_981) begin
          ways_3_metas_76_mru <= 1'b0;
        end
        if(_zz_982) begin
          ways_3_metas_77_mru <= 1'b0;
        end
        if(_zz_983) begin
          ways_3_metas_78_mru <= 1'b0;
        end
        if(_zz_984) begin
          ways_3_metas_79_mru <= 1'b0;
        end
        if(_zz_985) begin
          ways_3_metas_80_mru <= 1'b0;
        end
        if(_zz_986) begin
          ways_3_metas_81_mru <= 1'b0;
        end
        if(_zz_987) begin
          ways_3_metas_82_mru <= 1'b0;
        end
        if(_zz_988) begin
          ways_3_metas_83_mru <= 1'b0;
        end
        if(_zz_989) begin
          ways_3_metas_84_mru <= 1'b0;
        end
        if(_zz_990) begin
          ways_3_metas_85_mru <= 1'b0;
        end
        if(_zz_991) begin
          ways_3_metas_86_mru <= 1'b0;
        end
        if(_zz_992) begin
          ways_3_metas_87_mru <= 1'b0;
        end
        if(_zz_993) begin
          ways_3_metas_88_mru <= 1'b0;
        end
        if(_zz_994) begin
          ways_3_metas_89_mru <= 1'b0;
        end
        if(_zz_995) begin
          ways_3_metas_90_mru <= 1'b0;
        end
        if(_zz_996) begin
          ways_3_metas_91_mru <= 1'b0;
        end
        if(_zz_997) begin
          ways_3_metas_92_mru <= 1'b0;
        end
        if(_zz_998) begin
          ways_3_metas_93_mru <= 1'b0;
        end
        if(_zz_999) begin
          ways_3_metas_94_mru <= 1'b0;
        end
        if(_zz_1000) begin
          ways_3_metas_95_mru <= 1'b0;
        end
        if(_zz_1001) begin
          ways_3_metas_96_mru <= 1'b0;
        end
        if(_zz_1002) begin
          ways_3_metas_97_mru <= 1'b0;
        end
        if(_zz_1003) begin
          ways_3_metas_98_mru <= 1'b0;
        end
        if(_zz_1004) begin
          ways_3_metas_99_mru <= 1'b0;
        end
        if(_zz_1005) begin
          ways_3_metas_100_mru <= 1'b0;
        end
        if(_zz_1006) begin
          ways_3_metas_101_mru <= 1'b0;
        end
        if(_zz_1007) begin
          ways_3_metas_102_mru <= 1'b0;
        end
        if(_zz_1008) begin
          ways_3_metas_103_mru <= 1'b0;
        end
        if(_zz_1009) begin
          ways_3_metas_104_mru <= 1'b0;
        end
        if(_zz_1010) begin
          ways_3_metas_105_mru <= 1'b0;
        end
        if(_zz_1011) begin
          ways_3_metas_106_mru <= 1'b0;
        end
        if(_zz_1012) begin
          ways_3_metas_107_mru <= 1'b0;
        end
        if(_zz_1013) begin
          ways_3_metas_108_mru <= 1'b0;
        end
        if(_zz_1014) begin
          ways_3_metas_109_mru <= 1'b0;
        end
        if(_zz_1015) begin
          ways_3_metas_110_mru <= 1'b0;
        end
        if(_zz_1016) begin
          ways_3_metas_111_mru <= 1'b0;
        end
        if(_zz_1017) begin
          ways_3_metas_112_mru <= 1'b0;
        end
        if(_zz_1018) begin
          ways_3_metas_113_mru <= 1'b0;
        end
        if(_zz_1019) begin
          ways_3_metas_114_mru <= 1'b0;
        end
        if(_zz_1020) begin
          ways_3_metas_115_mru <= 1'b0;
        end
        if(_zz_1021) begin
          ways_3_metas_116_mru <= 1'b0;
        end
        if(_zz_1022) begin
          ways_3_metas_117_mru <= 1'b0;
        end
        if(_zz_1023) begin
          ways_3_metas_118_mru <= 1'b0;
        end
        if(_zz_1024) begin
          ways_3_metas_119_mru <= 1'b0;
        end
        if(_zz_1025) begin
          ways_3_metas_120_mru <= 1'b0;
        end
        if(_zz_1026) begin
          ways_3_metas_121_mru <= 1'b0;
        end
        if(_zz_1027) begin
          ways_3_metas_122_mru <= 1'b0;
        end
        if(_zz_1028) begin
          ways_3_metas_123_mru <= 1'b0;
        end
        if(_zz_1029) begin
          ways_3_metas_124_mru <= 1'b0;
        end
        if(_zz_1030) begin
          ways_3_metas_125_mru <= 1'b0;
        end
        if(_zz_1031) begin
          ways_3_metas_126_mru <= 1'b0;
        end
        if(_zz_1032) begin
          ways_3_metas_127_mru <= 1'b0;
        end
        if(_zz_905) begin
          ways_3_metas_0_vld <= 1'b0;
        end
        if(_zz_906) begin
          ways_3_metas_1_vld <= 1'b0;
        end
        if(_zz_907) begin
          ways_3_metas_2_vld <= 1'b0;
        end
        if(_zz_908) begin
          ways_3_metas_3_vld <= 1'b0;
        end
        if(_zz_909) begin
          ways_3_metas_4_vld <= 1'b0;
        end
        if(_zz_910) begin
          ways_3_metas_5_vld <= 1'b0;
        end
        if(_zz_911) begin
          ways_3_metas_6_vld <= 1'b0;
        end
        if(_zz_912) begin
          ways_3_metas_7_vld <= 1'b0;
        end
        if(_zz_913) begin
          ways_3_metas_8_vld <= 1'b0;
        end
        if(_zz_914) begin
          ways_3_metas_9_vld <= 1'b0;
        end
        if(_zz_915) begin
          ways_3_metas_10_vld <= 1'b0;
        end
        if(_zz_916) begin
          ways_3_metas_11_vld <= 1'b0;
        end
        if(_zz_917) begin
          ways_3_metas_12_vld <= 1'b0;
        end
        if(_zz_918) begin
          ways_3_metas_13_vld <= 1'b0;
        end
        if(_zz_919) begin
          ways_3_metas_14_vld <= 1'b0;
        end
        if(_zz_920) begin
          ways_3_metas_15_vld <= 1'b0;
        end
        if(_zz_921) begin
          ways_3_metas_16_vld <= 1'b0;
        end
        if(_zz_922) begin
          ways_3_metas_17_vld <= 1'b0;
        end
        if(_zz_923) begin
          ways_3_metas_18_vld <= 1'b0;
        end
        if(_zz_924) begin
          ways_3_metas_19_vld <= 1'b0;
        end
        if(_zz_925) begin
          ways_3_metas_20_vld <= 1'b0;
        end
        if(_zz_926) begin
          ways_3_metas_21_vld <= 1'b0;
        end
        if(_zz_927) begin
          ways_3_metas_22_vld <= 1'b0;
        end
        if(_zz_928) begin
          ways_3_metas_23_vld <= 1'b0;
        end
        if(_zz_929) begin
          ways_3_metas_24_vld <= 1'b0;
        end
        if(_zz_930) begin
          ways_3_metas_25_vld <= 1'b0;
        end
        if(_zz_931) begin
          ways_3_metas_26_vld <= 1'b0;
        end
        if(_zz_932) begin
          ways_3_metas_27_vld <= 1'b0;
        end
        if(_zz_933) begin
          ways_3_metas_28_vld <= 1'b0;
        end
        if(_zz_934) begin
          ways_3_metas_29_vld <= 1'b0;
        end
        if(_zz_935) begin
          ways_3_metas_30_vld <= 1'b0;
        end
        if(_zz_936) begin
          ways_3_metas_31_vld <= 1'b0;
        end
        if(_zz_937) begin
          ways_3_metas_32_vld <= 1'b0;
        end
        if(_zz_938) begin
          ways_3_metas_33_vld <= 1'b0;
        end
        if(_zz_939) begin
          ways_3_metas_34_vld <= 1'b0;
        end
        if(_zz_940) begin
          ways_3_metas_35_vld <= 1'b0;
        end
        if(_zz_941) begin
          ways_3_metas_36_vld <= 1'b0;
        end
        if(_zz_942) begin
          ways_3_metas_37_vld <= 1'b0;
        end
        if(_zz_943) begin
          ways_3_metas_38_vld <= 1'b0;
        end
        if(_zz_944) begin
          ways_3_metas_39_vld <= 1'b0;
        end
        if(_zz_945) begin
          ways_3_metas_40_vld <= 1'b0;
        end
        if(_zz_946) begin
          ways_3_metas_41_vld <= 1'b0;
        end
        if(_zz_947) begin
          ways_3_metas_42_vld <= 1'b0;
        end
        if(_zz_948) begin
          ways_3_metas_43_vld <= 1'b0;
        end
        if(_zz_949) begin
          ways_3_metas_44_vld <= 1'b0;
        end
        if(_zz_950) begin
          ways_3_metas_45_vld <= 1'b0;
        end
        if(_zz_951) begin
          ways_3_metas_46_vld <= 1'b0;
        end
        if(_zz_952) begin
          ways_3_metas_47_vld <= 1'b0;
        end
        if(_zz_953) begin
          ways_3_metas_48_vld <= 1'b0;
        end
        if(_zz_954) begin
          ways_3_metas_49_vld <= 1'b0;
        end
        if(_zz_955) begin
          ways_3_metas_50_vld <= 1'b0;
        end
        if(_zz_956) begin
          ways_3_metas_51_vld <= 1'b0;
        end
        if(_zz_957) begin
          ways_3_metas_52_vld <= 1'b0;
        end
        if(_zz_958) begin
          ways_3_metas_53_vld <= 1'b0;
        end
        if(_zz_959) begin
          ways_3_metas_54_vld <= 1'b0;
        end
        if(_zz_960) begin
          ways_3_metas_55_vld <= 1'b0;
        end
        if(_zz_961) begin
          ways_3_metas_56_vld <= 1'b0;
        end
        if(_zz_962) begin
          ways_3_metas_57_vld <= 1'b0;
        end
        if(_zz_963) begin
          ways_3_metas_58_vld <= 1'b0;
        end
        if(_zz_964) begin
          ways_3_metas_59_vld <= 1'b0;
        end
        if(_zz_965) begin
          ways_3_metas_60_vld <= 1'b0;
        end
        if(_zz_966) begin
          ways_3_metas_61_vld <= 1'b0;
        end
        if(_zz_967) begin
          ways_3_metas_62_vld <= 1'b0;
        end
        if(_zz_968) begin
          ways_3_metas_63_vld <= 1'b0;
        end
        if(_zz_969) begin
          ways_3_metas_64_vld <= 1'b0;
        end
        if(_zz_970) begin
          ways_3_metas_65_vld <= 1'b0;
        end
        if(_zz_971) begin
          ways_3_metas_66_vld <= 1'b0;
        end
        if(_zz_972) begin
          ways_3_metas_67_vld <= 1'b0;
        end
        if(_zz_973) begin
          ways_3_metas_68_vld <= 1'b0;
        end
        if(_zz_974) begin
          ways_3_metas_69_vld <= 1'b0;
        end
        if(_zz_975) begin
          ways_3_metas_70_vld <= 1'b0;
        end
        if(_zz_976) begin
          ways_3_metas_71_vld <= 1'b0;
        end
        if(_zz_977) begin
          ways_3_metas_72_vld <= 1'b0;
        end
        if(_zz_978) begin
          ways_3_metas_73_vld <= 1'b0;
        end
        if(_zz_979) begin
          ways_3_metas_74_vld <= 1'b0;
        end
        if(_zz_980) begin
          ways_3_metas_75_vld <= 1'b0;
        end
        if(_zz_981) begin
          ways_3_metas_76_vld <= 1'b0;
        end
        if(_zz_982) begin
          ways_3_metas_77_vld <= 1'b0;
        end
        if(_zz_983) begin
          ways_3_metas_78_vld <= 1'b0;
        end
        if(_zz_984) begin
          ways_3_metas_79_vld <= 1'b0;
        end
        if(_zz_985) begin
          ways_3_metas_80_vld <= 1'b0;
        end
        if(_zz_986) begin
          ways_3_metas_81_vld <= 1'b0;
        end
        if(_zz_987) begin
          ways_3_metas_82_vld <= 1'b0;
        end
        if(_zz_988) begin
          ways_3_metas_83_vld <= 1'b0;
        end
        if(_zz_989) begin
          ways_3_metas_84_vld <= 1'b0;
        end
        if(_zz_990) begin
          ways_3_metas_85_vld <= 1'b0;
        end
        if(_zz_991) begin
          ways_3_metas_86_vld <= 1'b0;
        end
        if(_zz_992) begin
          ways_3_metas_87_vld <= 1'b0;
        end
        if(_zz_993) begin
          ways_3_metas_88_vld <= 1'b0;
        end
        if(_zz_994) begin
          ways_3_metas_89_vld <= 1'b0;
        end
        if(_zz_995) begin
          ways_3_metas_90_vld <= 1'b0;
        end
        if(_zz_996) begin
          ways_3_metas_91_vld <= 1'b0;
        end
        if(_zz_997) begin
          ways_3_metas_92_vld <= 1'b0;
        end
        if(_zz_998) begin
          ways_3_metas_93_vld <= 1'b0;
        end
        if(_zz_999) begin
          ways_3_metas_94_vld <= 1'b0;
        end
        if(_zz_1000) begin
          ways_3_metas_95_vld <= 1'b0;
        end
        if(_zz_1001) begin
          ways_3_metas_96_vld <= 1'b0;
        end
        if(_zz_1002) begin
          ways_3_metas_97_vld <= 1'b0;
        end
        if(_zz_1003) begin
          ways_3_metas_98_vld <= 1'b0;
        end
        if(_zz_1004) begin
          ways_3_metas_99_vld <= 1'b0;
        end
        if(_zz_1005) begin
          ways_3_metas_100_vld <= 1'b0;
        end
        if(_zz_1006) begin
          ways_3_metas_101_vld <= 1'b0;
        end
        if(_zz_1007) begin
          ways_3_metas_102_vld <= 1'b0;
        end
        if(_zz_1008) begin
          ways_3_metas_103_vld <= 1'b0;
        end
        if(_zz_1009) begin
          ways_3_metas_104_vld <= 1'b0;
        end
        if(_zz_1010) begin
          ways_3_metas_105_vld <= 1'b0;
        end
        if(_zz_1011) begin
          ways_3_metas_106_vld <= 1'b0;
        end
        if(_zz_1012) begin
          ways_3_metas_107_vld <= 1'b0;
        end
        if(_zz_1013) begin
          ways_3_metas_108_vld <= 1'b0;
        end
        if(_zz_1014) begin
          ways_3_metas_109_vld <= 1'b0;
        end
        if(_zz_1015) begin
          ways_3_metas_110_vld <= 1'b0;
        end
        if(_zz_1016) begin
          ways_3_metas_111_vld <= 1'b0;
        end
        if(_zz_1017) begin
          ways_3_metas_112_vld <= 1'b0;
        end
        if(_zz_1018) begin
          ways_3_metas_113_vld <= 1'b0;
        end
        if(_zz_1019) begin
          ways_3_metas_114_vld <= 1'b0;
        end
        if(_zz_1020) begin
          ways_3_metas_115_vld <= 1'b0;
        end
        if(_zz_1021) begin
          ways_3_metas_116_vld <= 1'b0;
        end
        if(_zz_1022) begin
          ways_3_metas_117_vld <= 1'b0;
        end
        if(_zz_1023) begin
          ways_3_metas_118_vld <= 1'b0;
        end
        if(_zz_1024) begin
          ways_3_metas_119_vld <= 1'b0;
        end
        if(_zz_1025) begin
          ways_3_metas_120_vld <= 1'b0;
        end
        if(_zz_1026) begin
          ways_3_metas_121_vld <= 1'b0;
        end
        if(_zz_1027) begin
          ways_3_metas_122_vld <= 1'b0;
        end
        if(_zz_1028) begin
          ways_3_metas_123_vld <= 1'b0;
        end
        if(_zz_1029) begin
          ways_3_metas_124_vld <= 1'b0;
        end
        if(_zz_1030) begin
          ways_3_metas_125_vld <= 1'b0;
        end
        if(_zz_1031) begin
          ways_3_metas_126_vld <= 1'b0;
        end
        if(_zz_1032) begin
          ways_3_metas_127_vld <= 1'b0;
        end
      end else begin
        if(when_DCache_l217_3) begin
          if(cache_hit_3) begin
            if(_zz_776) begin
              ways_3_metas_0_mru <= 1'b1;
            end
            if(_zz_777) begin
              ways_3_metas_1_mru <= 1'b1;
            end
            if(_zz_778) begin
              ways_3_metas_2_mru <= 1'b1;
            end
            if(_zz_779) begin
              ways_3_metas_3_mru <= 1'b1;
            end
            if(_zz_780) begin
              ways_3_metas_4_mru <= 1'b1;
            end
            if(_zz_781) begin
              ways_3_metas_5_mru <= 1'b1;
            end
            if(_zz_782) begin
              ways_3_metas_6_mru <= 1'b1;
            end
            if(_zz_783) begin
              ways_3_metas_7_mru <= 1'b1;
            end
            if(_zz_784) begin
              ways_3_metas_8_mru <= 1'b1;
            end
            if(_zz_785) begin
              ways_3_metas_9_mru <= 1'b1;
            end
            if(_zz_786) begin
              ways_3_metas_10_mru <= 1'b1;
            end
            if(_zz_787) begin
              ways_3_metas_11_mru <= 1'b1;
            end
            if(_zz_788) begin
              ways_3_metas_12_mru <= 1'b1;
            end
            if(_zz_789) begin
              ways_3_metas_13_mru <= 1'b1;
            end
            if(_zz_790) begin
              ways_3_metas_14_mru <= 1'b1;
            end
            if(_zz_791) begin
              ways_3_metas_15_mru <= 1'b1;
            end
            if(_zz_792) begin
              ways_3_metas_16_mru <= 1'b1;
            end
            if(_zz_793) begin
              ways_3_metas_17_mru <= 1'b1;
            end
            if(_zz_794) begin
              ways_3_metas_18_mru <= 1'b1;
            end
            if(_zz_795) begin
              ways_3_metas_19_mru <= 1'b1;
            end
            if(_zz_796) begin
              ways_3_metas_20_mru <= 1'b1;
            end
            if(_zz_797) begin
              ways_3_metas_21_mru <= 1'b1;
            end
            if(_zz_798) begin
              ways_3_metas_22_mru <= 1'b1;
            end
            if(_zz_799) begin
              ways_3_metas_23_mru <= 1'b1;
            end
            if(_zz_800) begin
              ways_3_metas_24_mru <= 1'b1;
            end
            if(_zz_801) begin
              ways_3_metas_25_mru <= 1'b1;
            end
            if(_zz_802) begin
              ways_3_metas_26_mru <= 1'b1;
            end
            if(_zz_803) begin
              ways_3_metas_27_mru <= 1'b1;
            end
            if(_zz_804) begin
              ways_3_metas_28_mru <= 1'b1;
            end
            if(_zz_805) begin
              ways_3_metas_29_mru <= 1'b1;
            end
            if(_zz_806) begin
              ways_3_metas_30_mru <= 1'b1;
            end
            if(_zz_807) begin
              ways_3_metas_31_mru <= 1'b1;
            end
            if(_zz_808) begin
              ways_3_metas_32_mru <= 1'b1;
            end
            if(_zz_809) begin
              ways_3_metas_33_mru <= 1'b1;
            end
            if(_zz_810) begin
              ways_3_metas_34_mru <= 1'b1;
            end
            if(_zz_811) begin
              ways_3_metas_35_mru <= 1'b1;
            end
            if(_zz_812) begin
              ways_3_metas_36_mru <= 1'b1;
            end
            if(_zz_813) begin
              ways_3_metas_37_mru <= 1'b1;
            end
            if(_zz_814) begin
              ways_3_metas_38_mru <= 1'b1;
            end
            if(_zz_815) begin
              ways_3_metas_39_mru <= 1'b1;
            end
            if(_zz_816) begin
              ways_3_metas_40_mru <= 1'b1;
            end
            if(_zz_817) begin
              ways_3_metas_41_mru <= 1'b1;
            end
            if(_zz_818) begin
              ways_3_metas_42_mru <= 1'b1;
            end
            if(_zz_819) begin
              ways_3_metas_43_mru <= 1'b1;
            end
            if(_zz_820) begin
              ways_3_metas_44_mru <= 1'b1;
            end
            if(_zz_821) begin
              ways_3_metas_45_mru <= 1'b1;
            end
            if(_zz_822) begin
              ways_3_metas_46_mru <= 1'b1;
            end
            if(_zz_823) begin
              ways_3_metas_47_mru <= 1'b1;
            end
            if(_zz_824) begin
              ways_3_metas_48_mru <= 1'b1;
            end
            if(_zz_825) begin
              ways_3_metas_49_mru <= 1'b1;
            end
            if(_zz_826) begin
              ways_3_metas_50_mru <= 1'b1;
            end
            if(_zz_827) begin
              ways_3_metas_51_mru <= 1'b1;
            end
            if(_zz_828) begin
              ways_3_metas_52_mru <= 1'b1;
            end
            if(_zz_829) begin
              ways_3_metas_53_mru <= 1'b1;
            end
            if(_zz_830) begin
              ways_3_metas_54_mru <= 1'b1;
            end
            if(_zz_831) begin
              ways_3_metas_55_mru <= 1'b1;
            end
            if(_zz_832) begin
              ways_3_metas_56_mru <= 1'b1;
            end
            if(_zz_833) begin
              ways_3_metas_57_mru <= 1'b1;
            end
            if(_zz_834) begin
              ways_3_metas_58_mru <= 1'b1;
            end
            if(_zz_835) begin
              ways_3_metas_59_mru <= 1'b1;
            end
            if(_zz_836) begin
              ways_3_metas_60_mru <= 1'b1;
            end
            if(_zz_837) begin
              ways_3_metas_61_mru <= 1'b1;
            end
            if(_zz_838) begin
              ways_3_metas_62_mru <= 1'b1;
            end
            if(_zz_839) begin
              ways_3_metas_63_mru <= 1'b1;
            end
            if(_zz_840) begin
              ways_3_metas_64_mru <= 1'b1;
            end
            if(_zz_841) begin
              ways_3_metas_65_mru <= 1'b1;
            end
            if(_zz_842) begin
              ways_3_metas_66_mru <= 1'b1;
            end
            if(_zz_843) begin
              ways_3_metas_67_mru <= 1'b1;
            end
            if(_zz_844) begin
              ways_3_metas_68_mru <= 1'b1;
            end
            if(_zz_845) begin
              ways_3_metas_69_mru <= 1'b1;
            end
            if(_zz_846) begin
              ways_3_metas_70_mru <= 1'b1;
            end
            if(_zz_847) begin
              ways_3_metas_71_mru <= 1'b1;
            end
            if(_zz_848) begin
              ways_3_metas_72_mru <= 1'b1;
            end
            if(_zz_849) begin
              ways_3_metas_73_mru <= 1'b1;
            end
            if(_zz_850) begin
              ways_3_metas_74_mru <= 1'b1;
            end
            if(_zz_851) begin
              ways_3_metas_75_mru <= 1'b1;
            end
            if(_zz_852) begin
              ways_3_metas_76_mru <= 1'b1;
            end
            if(_zz_853) begin
              ways_3_metas_77_mru <= 1'b1;
            end
            if(_zz_854) begin
              ways_3_metas_78_mru <= 1'b1;
            end
            if(_zz_855) begin
              ways_3_metas_79_mru <= 1'b1;
            end
            if(_zz_856) begin
              ways_3_metas_80_mru <= 1'b1;
            end
            if(_zz_857) begin
              ways_3_metas_81_mru <= 1'b1;
            end
            if(_zz_858) begin
              ways_3_metas_82_mru <= 1'b1;
            end
            if(_zz_859) begin
              ways_3_metas_83_mru <= 1'b1;
            end
            if(_zz_860) begin
              ways_3_metas_84_mru <= 1'b1;
            end
            if(_zz_861) begin
              ways_3_metas_85_mru <= 1'b1;
            end
            if(_zz_862) begin
              ways_3_metas_86_mru <= 1'b1;
            end
            if(_zz_863) begin
              ways_3_metas_87_mru <= 1'b1;
            end
            if(_zz_864) begin
              ways_3_metas_88_mru <= 1'b1;
            end
            if(_zz_865) begin
              ways_3_metas_89_mru <= 1'b1;
            end
            if(_zz_866) begin
              ways_3_metas_90_mru <= 1'b1;
            end
            if(_zz_867) begin
              ways_3_metas_91_mru <= 1'b1;
            end
            if(_zz_868) begin
              ways_3_metas_92_mru <= 1'b1;
            end
            if(_zz_869) begin
              ways_3_metas_93_mru <= 1'b1;
            end
            if(_zz_870) begin
              ways_3_metas_94_mru <= 1'b1;
            end
            if(_zz_871) begin
              ways_3_metas_95_mru <= 1'b1;
            end
            if(_zz_872) begin
              ways_3_metas_96_mru <= 1'b1;
            end
            if(_zz_873) begin
              ways_3_metas_97_mru <= 1'b1;
            end
            if(_zz_874) begin
              ways_3_metas_98_mru <= 1'b1;
            end
            if(_zz_875) begin
              ways_3_metas_99_mru <= 1'b1;
            end
            if(_zz_876) begin
              ways_3_metas_100_mru <= 1'b1;
            end
            if(_zz_877) begin
              ways_3_metas_101_mru <= 1'b1;
            end
            if(_zz_878) begin
              ways_3_metas_102_mru <= 1'b1;
            end
            if(_zz_879) begin
              ways_3_metas_103_mru <= 1'b1;
            end
            if(_zz_880) begin
              ways_3_metas_104_mru <= 1'b1;
            end
            if(_zz_881) begin
              ways_3_metas_105_mru <= 1'b1;
            end
            if(_zz_882) begin
              ways_3_metas_106_mru <= 1'b1;
            end
            if(_zz_883) begin
              ways_3_metas_107_mru <= 1'b1;
            end
            if(_zz_884) begin
              ways_3_metas_108_mru <= 1'b1;
            end
            if(_zz_885) begin
              ways_3_metas_109_mru <= 1'b1;
            end
            if(_zz_886) begin
              ways_3_metas_110_mru <= 1'b1;
            end
            if(_zz_887) begin
              ways_3_metas_111_mru <= 1'b1;
            end
            if(_zz_888) begin
              ways_3_metas_112_mru <= 1'b1;
            end
            if(_zz_889) begin
              ways_3_metas_113_mru <= 1'b1;
            end
            if(_zz_890) begin
              ways_3_metas_114_mru <= 1'b1;
            end
            if(_zz_891) begin
              ways_3_metas_115_mru <= 1'b1;
            end
            if(_zz_892) begin
              ways_3_metas_116_mru <= 1'b1;
            end
            if(_zz_893) begin
              ways_3_metas_117_mru <= 1'b1;
            end
            if(_zz_894) begin
              ways_3_metas_118_mru <= 1'b1;
            end
            if(_zz_895) begin
              ways_3_metas_119_mru <= 1'b1;
            end
            if(_zz_896) begin
              ways_3_metas_120_mru <= 1'b1;
            end
            if(_zz_897) begin
              ways_3_metas_121_mru <= 1'b1;
            end
            if(_zz_898) begin
              ways_3_metas_122_mru <= 1'b1;
            end
            if(_zz_899) begin
              ways_3_metas_123_mru <= 1'b1;
            end
            if(_zz_900) begin
              ways_3_metas_124_mru <= 1'b1;
            end
            if(_zz_901) begin
              ways_3_metas_125_mru <= 1'b1;
            end
            if(_zz_902) begin
              ways_3_metas_126_mru <= 1'b1;
            end
            if(_zz_903) begin
              ways_3_metas_127_mru <= 1'b1;
            end
          end else begin
            if(_zz_776) begin
              ways_3_metas_0_mru <= 1'b0;
            end
            if(_zz_777) begin
              ways_3_metas_1_mru <= 1'b0;
            end
            if(_zz_778) begin
              ways_3_metas_2_mru <= 1'b0;
            end
            if(_zz_779) begin
              ways_3_metas_3_mru <= 1'b0;
            end
            if(_zz_780) begin
              ways_3_metas_4_mru <= 1'b0;
            end
            if(_zz_781) begin
              ways_3_metas_5_mru <= 1'b0;
            end
            if(_zz_782) begin
              ways_3_metas_6_mru <= 1'b0;
            end
            if(_zz_783) begin
              ways_3_metas_7_mru <= 1'b0;
            end
            if(_zz_784) begin
              ways_3_metas_8_mru <= 1'b0;
            end
            if(_zz_785) begin
              ways_3_metas_9_mru <= 1'b0;
            end
            if(_zz_786) begin
              ways_3_metas_10_mru <= 1'b0;
            end
            if(_zz_787) begin
              ways_3_metas_11_mru <= 1'b0;
            end
            if(_zz_788) begin
              ways_3_metas_12_mru <= 1'b0;
            end
            if(_zz_789) begin
              ways_3_metas_13_mru <= 1'b0;
            end
            if(_zz_790) begin
              ways_3_metas_14_mru <= 1'b0;
            end
            if(_zz_791) begin
              ways_3_metas_15_mru <= 1'b0;
            end
            if(_zz_792) begin
              ways_3_metas_16_mru <= 1'b0;
            end
            if(_zz_793) begin
              ways_3_metas_17_mru <= 1'b0;
            end
            if(_zz_794) begin
              ways_3_metas_18_mru <= 1'b0;
            end
            if(_zz_795) begin
              ways_3_metas_19_mru <= 1'b0;
            end
            if(_zz_796) begin
              ways_3_metas_20_mru <= 1'b0;
            end
            if(_zz_797) begin
              ways_3_metas_21_mru <= 1'b0;
            end
            if(_zz_798) begin
              ways_3_metas_22_mru <= 1'b0;
            end
            if(_zz_799) begin
              ways_3_metas_23_mru <= 1'b0;
            end
            if(_zz_800) begin
              ways_3_metas_24_mru <= 1'b0;
            end
            if(_zz_801) begin
              ways_3_metas_25_mru <= 1'b0;
            end
            if(_zz_802) begin
              ways_3_metas_26_mru <= 1'b0;
            end
            if(_zz_803) begin
              ways_3_metas_27_mru <= 1'b0;
            end
            if(_zz_804) begin
              ways_3_metas_28_mru <= 1'b0;
            end
            if(_zz_805) begin
              ways_3_metas_29_mru <= 1'b0;
            end
            if(_zz_806) begin
              ways_3_metas_30_mru <= 1'b0;
            end
            if(_zz_807) begin
              ways_3_metas_31_mru <= 1'b0;
            end
            if(_zz_808) begin
              ways_3_metas_32_mru <= 1'b0;
            end
            if(_zz_809) begin
              ways_3_metas_33_mru <= 1'b0;
            end
            if(_zz_810) begin
              ways_3_metas_34_mru <= 1'b0;
            end
            if(_zz_811) begin
              ways_3_metas_35_mru <= 1'b0;
            end
            if(_zz_812) begin
              ways_3_metas_36_mru <= 1'b0;
            end
            if(_zz_813) begin
              ways_3_metas_37_mru <= 1'b0;
            end
            if(_zz_814) begin
              ways_3_metas_38_mru <= 1'b0;
            end
            if(_zz_815) begin
              ways_3_metas_39_mru <= 1'b0;
            end
            if(_zz_816) begin
              ways_3_metas_40_mru <= 1'b0;
            end
            if(_zz_817) begin
              ways_3_metas_41_mru <= 1'b0;
            end
            if(_zz_818) begin
              ways_3_metas_42_mru <= 1'b0;
            end
            if(_zz_819) begin
              ways_3_metas_43_mru <= 1'b0;
            end
            if(_zz_820) begin
              ways_3_metas_44_mru <= 1'b0;
            end
            if(_zz_821) begin
              ways_3_metas_45_mru <= 1'b0;
            end
            if(_zz_822) begin
              ways_3_metas_46_mru <= 1'b0;
            end
            if(_zz_823) begin
              ways_3_metas_47_mru <= 1'b0;
            end
            if(_zz_824) begin
              ways_3_metas_48_mru <= 1'b0;
            end
            if(_zz_825) begin
              ways_3_metas_49_mru <= 1'b0;
            end
            if(_zz_826) begin
              ways_3_metas_50_mru <= 1'b0;
            end
            if(_zz_827) begin
              ways_3_metas_51_mru <= 1'b0;
            end
            if(_zz_828) begin
              ways_3_metas_52_mru <= 1'b0;
            end
            if(_zz_829) begin
              ways_3_metas_53_mru <= 1'b0;
            end
            if(_zz_830) begin
              ways_3_metas_54_mru <= 1'b0;
            end
            if(_zz_831) begin
              ways_3_metas_55_mru <= 1'b0;
            end
            if(_zz_832) begin
              ways_3_metas_56_mru <= 1'b0;
            end
            if(_zz_833) begin
              ways_3_metas_57_mru <= 1'b0;
            end
            if(_zz_834) begin
              ways_3_metas_58_mru <= 1'b0;
            end
            if(_zz_835) begin
              ways_3_metas_59_mru <= 1'b0;
            end
            if(_zz_836) begin
              ways_3_metas_60_mru <= 1'b0;
            end
            if(_zz_837) begin
              ways_3_metas_61_mru <= 1'b0;
            end
            if(_zz_838) begin
              ways_3_metas_62_mru <= 1'b0;
            end
            if(_zz_839) begin
              ways_3_metas_63_mru <= 1'b0;
            end
            if(_zz_840) begin
              ways_3_metas_64_mru <= 1'b0;
            end
            if(_zz_841) begin
              ways_3_metas_65_mru <= 1'b0;
            end
            if(_zz_842) begin
              ways_3_metas_66_mru <= 1'b0;
            end
            if(_zz_843) begin
              ways_3_metas_67_mru <= 1'b0;
            end
            if(_zz_844) begin
              ways_3_metas_68_mru <= 1'b0;
            end
            if(_zz_845) begin
              ways_3_metas_69_mru <= 1'b0;
            end
            if(_zz_846) begin
              ways_3_metas_70_mru <= 1'b0;
            end
            if(_zz_847) begin
              ways_3_metas_71_mru <= 1'b0;
            end
            if(_zz_848) begin
              ways_3_metas_72_mru <= 1'b0;
            end
            if(_zz_849) begin
              ways_3_metas_73_mru <= 1'b0;
            end
            if(_zz_850) begin
              ways_3_metas_74_mru <= 1'b0;
            end
            if(_zz_851) begin
              ways_3_metas_75_mru <= 1'b0;
            end
            if(_zz_852) begin
              ways_3_metas_76_mru <= 1'b0;
            end
            if(_zz_853) begin
              ways_3_metas_77_mru <= 1'b0;
            end
            if(_zz_854) begin
              ways_3_metas_78_mru <= 1'b0;
            end
            if(_zz_855) begin
              ways_3_metas_79_mru <= 1'b0;
            end
            if(_zz_856) begin
              ways_3_metas_80_mru <= 1'b0;
            end
            if(_zz_857) begin
              ways_3_metas_81_mru <= 1'b0;
            end
            if(_zz_858) begin
              ways_3_metas_82_mru <= 1'b0;
            end
            if(_zz_859) begin
              ways_3_metas_83_mru <= 1'b0;
            end
            if(_zz_860) begin
              ways_3_metas_84_mru <= 1'b0;
            end
            if(_zz_861) begin
              ways_3_metas_85_mru <= 1'b0;
            end
            if(_zz_862) begin
              ways_3_metas_86_mru <= 1'b0;
            end
            if(_zz_863) begin
              ways_3_metas_87_mru <= 1'b0;
            end
            if(_zz_864) begin
              ways_3_metas_88_mru <= 1'b0;
            end
            if(_zz_865) begin
              ways_3_metas_89_mru <= 1'b0;
            end
            if(_zz_866) begin
              ways_3_metas_90_mru <= 1'b0;
            end
            if(_zz_867) begin
              ways_3_metas_91_mru <= 1'b0;
            end
            if(_zz_868) begin
              ways_3_metas_92_mru <= 1'b0;
            end
            if(_zz_869) begin
              ways_3_metas_93_mru <= 1'b0;
            end
            if(_zz_870) begin
              ways_3_metas_94_mru <= 1'b0;
            end
            if(_zz_871) begin
              ways_3_metas_95_mru <= 1'b0;
            end
            if(_zz_872) begin
              ways_3_metas_96_mru <= 1'b0;
            end
            if(_zz_873) begin
              ways_3_metas_97_mru <= 1'b0;
            end
            if(_zz_874) begin
              ways_3_metas_98_mru <= 1'b0;
            end
            if(_zz_875) begin
              ways_3_metas_99_mru <= 1'b0;
            end
            if(_zz_876) begin
              ways_3_metas_100_mru <= 1'b0;
            end
            if(_zz_877) begin
              ways_3_metas_101_mru <= 1'b0;
            end
            if(_zz_878) begin
              ways_3_metas_102_mru <= 1'b0;
            end
            if(_zz_879) begin
              ways_3_metas_103_mru <= 1'b0;
            end
            if(_zz_880) begin
              ways_3_metas_104_mru <= 1'b0;
            end
            if(_zz_881) begin
              ways_3_metas_105_mru <= 1'b0;
            end
            if(_zz_882) begin
              ways_3_metas_106_mru <= 1'b0;
            end
            if(_zz_883) begin
              ways_3_metas_107_mru <= 1'b0;
            end
            if(_zz_884) begin
              ways_3_metas_108_mru <= 1'b0;
            end
            if(_zz_885) begin
              ways_3_metas_109_mru <= 1'b0;
            end
            if(_zz_886) begin
              ways_3_metas_110_mru <= 1'b0;
            end
            if(_zz_887) begin
              ways_3_metas_111_mru <= 1'b0;
            end
            if(_zz_888) begin
              ways_3_metas_112_mru <= 1'b0;
            end
            if(_zz_889) begin
              ways_3_metas_113_mru <= 1'b0;
            end
            if(_zz_890) begin
              ways_3_metas_114_mru <= 1'b0;
            end
            if(_zz_891) begin
              ways_3_metas_115_mru <= 1'b0;
            end
            if(_zz_892) begin
              ways_3_metas_116_mru <= 1'b0;
            end
            if(_zz_893) begin
              ways_3_metas_117_mru <= 1'b0;
            end
            if(_zz_894) begin
              ways_3_metas_118_mru <= 1'b0;
            end
            if(_zz_895) begin
              ways_3_metas_119_mru <= 1'b0;
            end
            if(_zz_896) begin
              ways_3_metas_120_mru <= 1'b0;
            end
            if(_zz_897) begin
              ways_3_metas_121_mru <= 1'b0;
            end
            if(_zz_898) begin
              ways_3_metas_122_mru <= 1'b0;
            end
            if(_zz_899) begin
              ways_3_metas_123_mru <= 1'b0;
            end
            if(_zz_900) begin
              ways_3_metas_124_mru <= 1'b0;
            end
            if(_zz_901) begin
              ways_3_metas_125_mru <= 1'b0;
            end
            if(_zz_902) begin
              ways_3_metas_126_mru <= 1'b0;
            end
            if(_zz_903) begin
              ways_3_metas_127_mru <= 1'b0;
            end
          end
        end else begin
          if(when_DCache_l224_3) begin
            if(_zz_776) begin
              ways_3_metas_0_mru <= 1'b1;
            end
            if(_zz_777) begin
              ways_3_metas_1_mru <= 1'b1;
            end
            if(_zz_778) begin
              ways_3_metas_2_mru <= 1'b1;
            end
            if(_zz_779) begin
              ways_3_metas_3_mru <= 1'b1;
            end
            if(_zz_780) begin
              ways_3_metas_4_mru <= 1'b1;
            end
            if(_zz_781) begin
              ways_3_metas_5_mru <= 1'b1;
            end
            if(_zz_782) begin
              ways_3_metas_6_mru <= 1'b1;
            end
            if(_zz_783) begin
              ways_3_metas_7_mru <= 1'b1;
            end
            if(_zz_784) begin
              ways_3_metas_8_mru <= 1'b1;
            end
            if(_zz_785) begin
              ways_3_metas_9_mru <= 1'b1;
            end
            if(_zz_786) begin
              ways_3_metas_10_mru <= 1'b1;
            end
            if(_zz_787) begin
              ways_3_metas_11_mru <= 1'b1;
            end
            if(_zz_788) begin
              ways_3_metas_12_mru <= 1'b1;
            end
            if(_zz_789) begin
              ways_3_metas_13_mru <= 1'b1;
            end
            if(_zz_790) begin
              ways_3_metas_14_mru <= 1'b1;
            end
            if(_zz_791) begin
              ways_3_metas_15_mru <= 1'b1;
            end
            if(_zz_792) begin
              ways_3_metas_16_mru <= 1'b1;
            end
            if(_zz_793) begin
              ways_3_metas_17_mru <= 1'b1;
            end
            if(_zz_794) begin
              ways_3_metas_18_mru <= 1'b1;
            end
            if(_zz_795) begin
              ways_3_metas_19_mru <= 1'b1;
            end
            if(_zz_796) begin
              ways_3_metas_20_mru <= 1'b1;
            end
            if(_zz_797) begin
              ways_3_metas_21_mru <= 1'b1;
            end
            if(_zz_798) begin
              ways_3_metas_22_mru <= 1'b1;
            end
            if(_zz_799) begin
              ways_3_metas_23_mru <= 1'b1;
            end
            if(_zz_800) begin
              ways_3_metas_24_mru <= 1'b1;
            end
            if(_zz_801) begin
              ways_3_metas_25_mru <= 1'b1;
            end
            if(_zz_802) begin
              ways_3_metas_26_mru <= 1'b1;
            end
            if(_zz_803) begin
              ways_3_metas_27_mru <= 1'b1;
            end
            if(_zz_804) begin
              ways_3_metas_28_mru <= 1'b1;
            end
            if(_zz_805) begin
              ways_3_metas_29_mru <= 1'b1;
            end
            if(_zz_806) begin
              ways_3_metas_30_mru <= 1'b1;
            end
            if(_zz_807) begin
              ways_3_metas_31_mru <= 1'b1;
            end
            if(_zz_808) begin
              ways_3_metas_32_mru <= 1'b1;
            end
            if(_zz_809) begin
              ways_3_metas_33_mru <= 1'b1;
            end
            if(_zz_810) begin
              ways_3_metas_34_mru <= 1'b1;
            end
            if(_zz_811) begin
              ways_3_metas_35_mru <= 1'b1;
            end
            if(_zz_812) begin
              ways_3_metas_36_mru <= 1'b1;
            end
            if(_zz_813) begin
              ways_3_metas_37_mru <= 1'b1;
            end
            if(_zz_814) begin
              ways_3_metas_38_mru <= 1'b1;
            end
            if(_zz_815) begin
              ways_3_metas_39_mru <= 1'b1;
            end
            if(_zz_816) begin
              ways_3_metas_40_mru <= 1'b1;
            end
            if(_zz_817) begin
              ways_3_metas_41_mru <= 1'b1;
            end
            if(_zz_818) begin
              ways_3_metas_42_mru <= 1'b1;
            end
            if(_zz_819) begin
              ways_3_metas_43_mru <= 1'b1;
            end
            if(_zz_820) begin
              ways_3_metas_44_mru <= 1'b1;
            end
            if(_zz_821) begin
              ways_3_metas_45_mru <= 1'b1;
            end
            if(_zz_822) begin
              ways_3_metas_46_mru <= 1'b1;
            end
            if(_zz_823) begin
              ways_3_metas_47_mru <= 1'b1;
            end
            if(_zz_824) begin
              ways_3_metas_48_mru <= 1'b1;
            end
            if(_zz_825) begin
              ways_3_metas_49_mru <= 1'b1;
            end
            if(_zz_826) begin
              ways_3_metas_50_mru <= 1'b1;
            end
            if(_zz_827) begin
              ways_3_metas_51_mru <= 1'b1;
            end
            if(_zz_828) begin
              ways_3_metas_52_mru <= 1'b1;
            end
            if(_zz_829) begin
              ways_3_metas_53_mru <= 1'b1;
            end
            if(_zz_830) begin
              ways_3_metas_54_mru <= 1'b1;
            end
            if(_zz_831) begin
              ways_3_metas_55_mru <= 1'b1;
            end
            if(_zz_832) begin
              ways_3_metas_56_mru <= 1'b1;
            end
            if(_zz_833) begin
              ways_3_metas_57_mru <= 1'b1;
            end
            if(_zz_834) begin
              ways_3_metas_58_mru <= 1'b1;
            end
            if(_zz_835) begin
              ways_3_metas_59_mru <= 1'b1;
            end
            if(_zz_836) begin
              ways_3_metas_60_mru <= 1'b1;
            end
            if(_zz_837) begin
              ways_3_metas_61_mru <= 1'b1;
            end
            if(_zz_838) begin
              ways_3_metas_62_mru <= 1'b1;
            end
            if(_zz_839) begin
              ways_3_metas_63_mru <= 1'b1;
            end
            if(_zz_840) begin
              ways_3_metas_64_mru <= 1'b1;
            end
            if(_zz_841) begin
              ways_3_metas_65_mru <= 1'b1;
            end
            if(_zz_842) begin
              ways_3_metas_66_mru <= 1'b1;
            end
            if(_zz_843) begin
              ways_3_metas_67_mru <= 1'b1;
            end
            if(_zz_844) begin
              ways_3_metas_68_mru <= 1'b1;
            end
            if(_zz_845) begin
              ways_3_metas_69_mru <= 1'b1;
            end
            if(_zz_846) begin
              ways_3_metas_70_mru <= 1'b1;
            end
            if(_zz_847) begin
              ways_3_metas_71_mru <= 1'b1;
            end
            if(_zz_848) begin
              ways_3_metas_72_mru <= 1'b1;
            end
            if(_zz_849) begin
              ways_3_metas_73_mru <= 1'b1;
            end
            if(_zz_850) begin
              ways_3_metas_74_mru <= 1'b1;
            end
            if(_zz_851) begin
              ways_3_metas_75_mru <= 1'b1;
            end
            if(_zz_852) begin
              ways_3_metas_76_mru <= 1'b1;
            end
            if(_zz_853) begin
              ways_3_metas_77_mru <= 1'b1;
            end
            if(_zz_854) begin
              ways_3_metas_78_mru <= 1'b1;
            end
            if(_zz_855) begin
              ways_3_metas_79_mru <= 1'b1;
            end
            if(_zz_856) begin
              ways_3_metas_80_mru <= 1'b1;
            end
            if(_zz_857) begin
              ways_3_metas_81_mru <= 1'b1;
            end
            if(_zz_858) begin
              ways_3_metas_82_mru <= 1'b1;
            end
            if(_zz_859) begin
              ways_3_metas_83_mru <= 1'b1;
            end
            if(_zz_860) begin
              ways_3_metas_84_mru <= 1'b1;
            end
            if(_zz_861) begin
              ways_3_metas_85_mru <= 1'b1;
            end
            if(_zz_862) begin
              ways_3_metas_86_mru <= 1'b1;
            end
            if(_zz_863) begin
              ways_3_metas_87_mru <= 1'b1;
            end
            if(_zz_864) begin
              ways_3_metas_88_mru <= 1'b1;
            end
            if(_zz_865) begin
              ways_3_metas_89_mru <= 1'b1;
            end
            if(_zz_866) begin
              ways_3_metas_90_mru <= 1'b1;
            end
            if(_zz_867) begin
              ways_3_metas_91_mru <= 1'b1;
            end
            if(_zz_868) begin
              ways_3_metas_92_mru <= 1'b1;
            end
            if(_zz_869) begin
              ways_3_metas_93_mru <= 1'b1;
            end
            if(_zz_870) begin
              ways_3_metas_94_mru <= 1'b1;
            end
            if(_zz_871) begin
              ways_3_metas_95_mru <= 1'b1;
            end
            if(_zz_872) begin
              ways_3_metas_96_mru <= 1'b1;
            end
            if(_zz_873) begin
              ways_3_metas_97_mru <= 1'b1;
            end
            if(_zz_874) begin
              ways_3_metas_98_mru <= 1'b1;
            end
            if(_zz_875) begin
              ways_3_metas_99_mru <= 1'b1;
            end
            if(_zz_876) begin
              ways_3_metas_100_mru <= 1'b1;
            end
            if(_zz_877) begin
              ways_3_metas_101_mru <= 1'b1;
            end
            if(_zz_878) begin
              ways_3_metas_102_mru <= 1'b1;
            end
            if(_zz_879) begin
              ways_3_metas_103_mru <= 1'b1;
            end
            if(_zz_880) begin
              ways_3_metas_104_mru <= 1'b1;
            end
            if(_zz_881) begin
              ways_3_metas_105_mru <= 1'b1;
            end
            if(_zz_882) begin
              ways_3_metas_106_mru <= 1'b1;
            end
            if(_zz_883) begin
              ways_3_metas_107_mru <= 1'b1;
            end
            if(_zz_884) begin
              ways_3_metas_108_mru <= 1'b1;
            end
            if(_zz_885) begin
              ways_3_metas_109_mru <= 1'b1;
            end
            if(_zz_886) begin
              ways_3_metas_110_mru <= 1'b1;
            end
            if(_zz_887) begin
              ways_3_metas_111_mru <= 1'b1;
            end
            if(_zz_888) begin
              ways_3_metas_112_mru <= 1'b1;
            end
            if(_zz_889) begin
              ways_3_metas_113_mru <= 1'b1;
            end
            if(_zz_890) begin
              ways_3_metas_114_mru <= 1'b1;
            end
            if(_zz_891) begin
              ways_3_metas_115_mru <= 1'b1;
            end
            if(_zz_892) begin
              ways_3_metas_116_mru <= 1'b1;
            end
            if(_zz_893) begin
              ways_3_metas_117_mru <= 1'b1;
            end
            if(_zz_894) begin
              ways_3_metas_118_mru <= 1'b1;
            end
            if(_zz_895) begin
              ways_3_metas_119_mru <= 1'b1;
            end
            if(_zz_896) begin
              ways_3_metas_120_mru <= 1'b1;
            end
            if(_zz_897) begin
              ways_3_metas_121_mru <= 1'b1;
            end
            if(_zz_898) begin
              ways_3_metas_122_mru <= 1'b1;
            end
            if(_zz_899) begin
              ways_3_metas_123_mru <= 1'b1;
            end
            if(_zz_900) begin
              ways_3_metas_124_mru <= 1'b1;
            end
            if(_zz_901) begin
              ways_3_metas_125_mru <= 1'b1;
            end
            if(_zz_902) begin
              ways_3_metas_126_mru <= 1'b1;
            end
            if(_zz_903) begin
              ways_3_metas_127_mru <= 1'b1;
            end
          end else begin
            if(when_DCache_l227_3) begin
              if(_zz_776) begin
                ways_3_metas_0_vld <= 1'b1;
              end
              if(_zz_777) begin
                ways_3_metas_1_vld <= 1'b1;
              end
              if(_zz_778) begin
                ways_3_metas_2_vld <= 1'b1;
              end
              if(_zz_779) begin
                ways_3_metas_3_vld <= 1'b1;
              end
              if(_zz_780) begin
                ways_3_metas_4_vld <= 1'b1;
              end
              if(_zz_781) begin
                ways_3_metas_5_vld <= 1'b1;
              end
              if(_zz_782) begin
                ways_3_metas_6_vld <= 1'b1;
              end
              if(_zz_783) begin
                ways_3_metas_7_vld <= 1'b1;
              end
              if(_zz_784) begin
                ways_3_metas_8_vld <= 1'b1;
              end
              if(_zz_785) begin
                ways_3_metas_9_vld <= 1'b1;
              end
              if(_zz_786) begin
                ways_3_metas_10_vld <= 1'b1;
              end
              if(_zz_787) begin
                ways_3_metas_11_vld <= 1'b1;
              end
              if(_zz_788) begin
                ways_3_metas_12_vld <= 1'b1;
              end
              if(_zz_789) begin
                ways_3_metas_13_vld <= 1'b1;
              end
              if(_zz_790) begin
                ways_3_metas_14_vld <= 1'b1;
              end
              if(_zz_791) begin
                ways_3_metas_15_vld <= 1'b1;
              end
              if(_zz_792) begin
                ways_3_metas_16_vld <= 1'b1;
              end
              if(_zz_793) begin
                ways_3_metas_17_vld <= 1'b1;
              end
              if(_zz_794) begin
                ways_3_metas_18_vld <= 1'b1;
              end
              if(_zz_795) begin
                ways_3_metas_19_vld <= 1'b1;
              end
              if(_zz_796) begin
                ways_3_metas_20_vld <= 1'b1;
              end
              if(_zz_797) begin
                ways_3_metas_21_vld <= 1'b1;
              end
              if(_zz_798) begin
                ways_3_metas_22_vld <= 1'b1;
              end
              if(_zz_799) begin
                ways_3_metas_23_vld <= 1'b1;
              end
              if(_zz_800) begin
                ways_3_metas_24_vld <= 1'b1;
              end
              if(_zz_801) begin
                ways_3_metas_25_vld <= 1'b1;
              end
              if(_zz_802) begin
                ways_3_metas_26_vld <= 1'b1;
              end
              if(_zz_803) begin
                ways_3_metas_27_vld <= 1'b1;
              end
              if(_zz_804) begin
                ways_3_metas_28_vld <= 1'b1;
              end
              if(_zz_805) begin
                ways_3_metas_29_vld <= 1'b1;
              end
              if(_zz_806) begin
                ways_3_metas_30_vld <= 1'b1;
              end
              if(_zz_807) begin
                ways_3_metas_31_vld <= 1'b1;
              end
              if(_zz_808) begin
                ways_3_metas_32_vld <= 1'b1;
              end
              if(_zz_809) begin
                ways_3_metas_33_vld <= 1'b1;
              end
              if(_zz_810) begin
                ways_3_metas_34_vld <= 1'b1;
              end
              if(_zz_811) begin
                ways_3_metas_35_vld <= 1'b1;
              end
              if(_zz_812) begin
                ways_3_metas_36_vld <= 1'b1;
              end
              if(_zz_813) begin
                ways_3_metas_37_vld <= 1'b1;
              end
              if(_zz_814) begin
                ways_3_metas_38_vld <= 1'b1;
              end
              if(_zz_815) begin
                ways_3_metas_39_vld <= 1'b1;
              end
              if(_zz_816) begin
                ways_3_metas_40_vld <= 1'b1;
              end
              if(_zz_817) begin
                ways_3_metas_41_vld <= 1'b1;
              end
              if(_zz_818) begin
                ways_3_metas_42_vld <= 1'b1;
              end
              if(_zz_819) begin
                ways_3_metas_43_vld <= 1'b1;
              end
              if(_zz_820) begin
                ways_3_metas_44_vld <= 1'b1;
              end
              if(_zz_821) begin
                ways_3_metas_45_vld <= 1'b1;
              end
              if(_zz_822) begin
                ways_3_metas_46_vld <= 1'b1;
              end
              if(_zz_823) begin
                ways_3_metas_47_vld <= 1'b1;
              end
              if(_zz_824) begin
                ways_3_metas_48_vld <= 1'b1;
              end
              if(_zz_825) begin
                ways_3_metas_49_vld <= 1'b1;
              end
              if(_zz_826) begin
                ways_3_metas_50_vld <= 1'b1;
              end
              if(_zz_827) begin
                ways_3_metas_51_vld <= 1'b1;
              end
              if(_zz_828) begin
                ways_3_metas_52_vld <= 1'b1;
              end
              if(_zz_829) begin
                ways_3_metas_53_vld <= 1'b1;
              end
              if(_zz_830) begin
                ways_3_metas_54_vld <= 1'b1;
              end
              if(_zz_831) begin
                ways_3_metas_55_vld <= 1'b1;
              end
              if(_zz_832) begin
                ways_3_metas_56_vld <= 1'b1;
              end
              if(_zz_833) begin
                ways_3_metas_57_vld <= 1'b1;
              end
              if(_zz_834) begin
                ways_3_metas_58_vld <= 1'b1;
              end
              if(_zz_835) begin
                ways_3_metas_59_vld <= 1'b1;
              end
              if(_zz_836) begin
                ways_3_metas_60_vld <= 1'b1;
              end
              if(_zz_837) begin
                ways_3_metas_61_vld <= 1'b1;
              end
              if(_zz_838) begin
                ways_3_metas_62_vld <= 1'b1;
              end
              if(_zz_839) begin
                ways_3_metas_63_vld <= 1'b1;
              end
              if(_zz_840) begin
                ways_3_metas_64_vld <= 1'b1;
              end
              if(_zz_841) begin
                ways_3_metas_65_vld <= 1'b1;
              end
              if(_zz_842) begin
                ways_3_metas_66_vld <= 1'b1;
              end
              if(_zz_843) begin
                ways_3_metas_67_vld <= 1'b1;
              end
              if(_zz_844) begin
                ways_3_metas_68_vld <= 1'b1;
              end
              if(_zz_845) begin
                ways_3_metas_69_vld <= 1'b1;
              end
              if(_zz_846) begin
                ways_3_metas_70_vld <= 1'b1;
              end
              if(_zz_847) begin
                ways_3_metas_71_vld <= 1'b1;
              end
              if(_zz_848) begin
                ways_3_metas_72_vld <= 1'b1;
              end
              if(_zz_849) begin
                ways_3_metas_73_vld <= 1'b1;
              end
              if(_zz_850) begin
                ways_3_metas_74_vld <= 1'b1;
              end
              if(_zz_851) begin
                ways_3_metas_75_vld <= 1'b1;
              end
              if(_zz_852) begin
                ways_3_metas_76_vld <= 1'b1;
              end
              if(_zz_853) begin
                ways_3_metas_77_vld <= 1'b1;
              end
              if(_zz_854) begin
                ways_3_metas_78_vld <= 1'b1;
              end
              if(_zz_855) begin
                ways_3_metas_79_vld <= 1'b1;
              end
              if(_zz_856) begin
                ways_3_metas_80_vld <= 1'b1;
              end
              if(_zz_857) begin
                ways_3_metas_81_vld <= 1'b1;
              end
              if(_zz_858) begin
                ways_3_metas_82_vld <= 1'b1;
              end
              if(_zz_859) begin
                ways_3_metas_83_vld <= 1'b1;
              end
              if(_zz_860) begin
                ways_3_metas_84_vld <= 1'b1;
              end
              if(_zz_861) begin
                ways_3_metas_85_vld <= 1'b1;
              end
              if(_zz_862) begin
                ways_3_metas_86_vld <= 1'b1;
              end
              if(_zz_863) begin
                ways_3_metas_87_vld <= 1'b1;
              end
              if(_zz_864) begin
                ways_3_metas_88_vld <= 1'b1;
              end
              if(_zz_865) begin
                ways_3_metas_89_vld <= 1'b1;
              end
              if(_zz_866) begin
                ways_3_metas_90_vld <= 1'b1;
              end
              if(_zz_867) begin
                ways_3_metas_91_vld <= 1'b1;
              end
              if(_zz_868) begin
                ways_3_metas_92_vld <= 1'b1;
              end
              if(_zz_869) begin
                ways_3_metas_93_vld <= 1'b1;
              end
              if(_zz_870) begin
                ways_3_metas_94_vld <= 1'b1;
              end
              if(_zz_871) begin
                ways_3_metas_95_vld <= 1'b1;
              end
              if(_zz_872) begin
                ways_3_metas_96_vld <= 1'b1;
              end
              if(_zz_873) begin
                ways_3_metas_97_vld <= 1'b1;
              end
              if(_zz_874) begin
                ways_3_metas_98_vld <= 1'b1;
              end
              if(_zz_875) begin
                ways_3_metas_99_vld <= 1'b1;
              end
              if(_zz_876) begin
                ways_3_metas_100_vld <= 1'b1;
              end
              if(_zz_877) begin
                ways_3_metas_101_vld <= 1'b1;
              end
              if(_zz_878) begin
                ways_3_metas_102_vld <= 1'b1;
              end
              if(_zz_879) begin
                ways_3_metas_103_vld <= 1'b1;
              end
              if(_zz_880) begin
                ways_3_metas_104_vld <= 1'b1;
              end
              if(_zz_881) begin
                ways_3_metas_105_vld <= 1'b1;
              end
              if(_zz_882) begin
                ways_3_metas_106_vld <= 1'b1;
              end
              if(_zz_883) begin
                ways_3_metas_107_vld <= 1'b1;
              end
              if(_zz_884) begin
                ways_3_metas_108_vld <= 1'b1;
              end
              if(_zz_885) begin
                ways_3_metas_109_vld <= 1'b1;
              end
              if(_zz_886) begin
                ways_3_metas_110_vld <= 1'b1;
              end
              if(_zz_887) begin
                ways_3_metas_111_vld <= 1'b1;
              end
              if(_zz_888) begin
                ways_3_metas_112_vld <= 1'b1;
              end
              if(_zz_889) begin
                ways_3_metas_113_vld <= 1'b1;
              end
              if(_zz_890) begin
                ways_3_metas_114_vld <= 1'b1;
              end
              if(_zz_891) begin
                ways_3_metas_115_vld <= 1'b1;
              end
              if(_zz_892) begin
                ways_3_metas_116_vld <= 1'b1;
              end
              if(_zz_893) begin
                ways_3_metas_117_vld <= 1'b1;
              end
              if(_zz_894) begin
                ways_3_metas_118_vld <= 1'b1;
              end
              if(_zz_895) begin
                ways_3_metas_119_vld <= 1'b1;
              end
              if(_zz_896) begin
                ways_3_metas_120_vld <= 1'b1;
              end
              if(_zz_897) begin
                ways_3_metas_121_vld <= 1'b1;
              end
              if(_zz_898) begin
                ways_3_metas_122_vld <= 1'b1;
              end
              if(_zz_899) begin
                ways_3_metas_123_vld <= 1'b1;
              end
              if(_zz_900) begin
                ways_3_metas_124_vld <= 1'b1;
              end
              if(_zz_901) begin
                ways_3_metas_125_vld <= 1'b1;
              end
              if(_zz_902) begin
                ways_3_metas_126_vld <= 1'b1;
              end
              if(_zz_903) begin
                ways_3_metas_127_vld <= 1'b1;
              end
            end
          end
        end
      end
      if(when_DCache_l232_3) begin
        if(_zz_776) begin
          ways_3_metas_0_tag <= cpu_tag;
        end
        if(_zz_777) begin
          ways_3_metas_1_tag <= cpu_tag;
        end
        if(_zz_778) begin
          ways_3_metas_2_tag <= cpu_tag;
        end
        if(_zz_779) begin
          ways_3_metas_3_tag <= cpu_tag;
        end
        if(_zz_780) begin
          ways_3_metas_4_tag <= cpu_tag;
        end
        if(_zz_781) begin
          ways_3_metas_5_tag <= cpu_tag;
        end
        if(_zz_782) begin
          ways_3_metas_6_tag <= cpu_tag;
        end
        if(_zz_783) begin
          ways_3_metas_7_tag <= cpu_tag;
        end
        if(_zz_784) begin
          ways_3_metas_8_tag <= cpu_tag;
        end
        if(_zz_785) begin
          ways_3_metas_9_tag <= cpu_tag;
        end
        if(_zz_786) begin
          ways_3_metas_10_tag <= cpu_tag;
        end
        if(_zz_787) begin
          ways_3_metas_11_tag <= cpu_tag;
        end
        if(_zz_788) begin
          ways_3_metas_12_tag <= cpu_tag;
        end
        if(_zz_789) begin
          ways_3_metas_13_tag <= cpu_tag;
        end
        if(_zz_790) begin
          ways_3_metas_14_tag <= cpu_tag;
        end
        if(_zz_791) begin
          ways_3_metas_15_tag <= cpu_tag;
        end
        if(_zz_792) begin
          ways_3_metas_16_tag <= cpu_tag;
        end
        if(_zz_793) begin
          ways_3_metas_17_tag <= cpu_tag;
        end
        if(_zz_794) begin
          ways_3_metas_18_tag <= cpu_tag;
        end
        if(_zz_795) begin
          ways_3_metas_19_tag <= cpu_tag;
        end
        if(_zz_796) begin
          ways_3_metas_20_tag <= cpu_tag;
        end
        if(_zz_797) begin
          ways_3_metas_21_tag <= cpu_tag;
        end
        if(_zz_798) begin
          ways_3_metas_22_tag <= cpu_tag;
        end
        if(_zz_799) begin
          ways_3_metas_23_tag <= cpu_tag;
        end
        if(_zz_800) begin
          ways_3_metas_24_tag <= cpu_tag;
        end
        if(_zz_801) begin
          ways_3_metas_25_tag <= cpu_tag;
        end
        if(_zz_802) begin
          ways_3_metas_26_tag <= cpu_tag;
        end
        if(_zz_803) begin
          ways_3_metas_27_tag <= cpu_tag;
        end
        if(_zz_804) begin
          ways_3_metas_28_tag <= cpu_tag;
        end
        if(_zz_805) begin
          ways_3_metas_29_tag <= cpu_tag;
        end
        if(_zz_806) begin
          ways_3_metas_30_tag <= cpu_tag;
        end
        if(_zz_807) begin
          ways_3_metas_31_tag <= cpu_tag;
        end
        if(_zz_808) begin
          ways_3_metas_32_tag <= cpu_tag;
        end
        if(_zz_809) begin
          ways_3_metas_33_tag <= cpu_tag;
        end
        if(_zz_810) begin
          ways_3_metas_34_tag <= cpu_tag;
        end
        if(_zz_811) begin
          ways_3_metas_35_tag <= cpu_tag;
        end
        if(_zz_812) begin
          ways_3_metas_36_tag <= cpu_tag;
        end
        if(_zz_813) begin
          ways_3_metas_37_tag <= cpu_tag;
        end
        if(_zz_814) begin
          ways_3_metas_38_tag <= cpu_tag;
        end
        if(_zz_815) begin
          ways_3_metas_39_tag <= cpu_tag;
        end
        if(_zz_816) begin
          ways_3_metas_40_tag <= cpu_tag;
        end
        if(_zz_817) begin
          ways_3_metas_41_tag <= cpu_tag;
        end
        if(_zz_818) begin
          ways_3_metas_42_tag <= cpu_tag;
        end
        if(_zz_819) begin
          ways_3_metas_43_tag <= cpu_tag;
        end
        if(_zz_820) begin
          ways_3_metas_44_tag <= cpu_tag;
        end
        if(_zz_821) begin
          ways_3_metas_45_tag <= cpu_tag;
        end
        if(_zz_822) begin
          ways_3_metas_46_tag <= cpu_tag;
        end
        if(_zz_823) begin
          ways_3_metas_47_tag <= cpu_tag;
        end
        if(_zz_824) begin
          ways_3_metas_48_tag <= cpu_tag;
        end
        if(_zz_825) begin
          ways_3_metas_49_tag <= cpu_tag;
        end
        if(_zz_826) begin
          ways_3_metas_50_tag <= cpu_tag;
        end
        if(_zz_827) begin
          ways_3_metas_51_tag <= cpu_tag;
        end
        if(_zz_828) begin
          ways_3_metas_52_tag <= cpu_tag;
        end
        if(_zz_829) begin
          ways_3_metas_53_tag <= cpu_tag;
        end
        if(_zz_830) begin
          ways_3_metas_54_tag <= cpu_tag;
        end
        if(_zz_831) begin
          ways_3_metas_55_tag <= cpu_tag;
        end
        if(_zz_832) begin
          ways_3_metas_56_tag <= cpu_tag;
        end
        if(_zz_833) begin
          ways_3_metas_57_tag <= cpu_tag;
        end
        if(_zz_834) begin
          ways_3_metas_58_tag <= cpu_tag;
        end
        if(_zz_835) begin
          ways_3_metas_59_tag <= cpu_tag;
        end
        if(_zz_836) begin
          ways_3_metas_60_tag <= cpu_tag;
        end
        if(_zz_837) begin
          ways_3_metas_61_tag <= cpu_tag;
        end
        if(_zz_838) begin
          ways_3_metas_62_tag <= cpu_tag;
        end
        if(_zz_839) begin
          ways_3_metas_63_tag <= cpu_tag;
        end
        if(_zz_840) begin
          ways_3_metas_64_tag <= cpu_tag;
        end
        if(_zz_841) begin
          ways_3_metas_65_tag <= cpu_tag;
        end
        if(_zz_842) begin
          ways_3_metas_66_tag <= cpu_tag;
        end
        if(_zz_843) begin
          ways_3_metas_67_tag <= cpu_tag;
        end
        if(_zz_844) begin
          ways_3_metas_68_tag <= cpu_tag;
        end
        if(_zz_845) begin
          ways_3_metas_69_tag <= cpu_tag;
        end
        if(_zz_846) begin
          ways_3_metas_70_tag <= cpu_tag;
        end
        if(_zz_847) begin
          ways_3_metas_71_tag <= cpu_tag;
        end
        if(_zz_848) begin
          ways_3_metas_72_tag <= cpu_tag;
        end
        if(_zz_849) begin
          ways_3_metas_73_tag <= cpu_tag;
        end
        if(_zz_850) begin
          ways_3_metas_74_tag <= cpu_tag;
        end
        if(_zz_851) begin
          ways_3_metas_75_tag <= cpu_tag;
        end
        if(_zz_852) begin
          ways_3_metas_76_tag <= cpu_tag;
        end
        if(_zz_853) begin
          ways_3_metas_77_tag <= cpu_tag;
        end
        if(_zz_854) begin
          ways_3_metas_78_tag <= cpu_tag;
        end
        if(_zz_855) begin
          ways_3_metas_79_tag <= cpu_tag;
        end
        if(_zz_856) begin
          ways_3_metas_80_tag <= cpu_tag;
        end
        if(_zz_857) begin
          ways_3_metas_81_tag <= cpu_tag;
        end
        if(_zz_858) begin
          ways_3_metas_82_tag <= cpu_tag;
        end
        if(_zz_859) begin
          ways_3_metas_83_tag <= cpu_tag;
        end
        if(_zz_860) begin
          ways_3_metas_84_tag <= cpu_tag;
        end
        if(_zz_861) begin
          ways_3_metas_85_tag <= cpu_tag;
        end
        if(_zz_862) begin
          ways_3_metas_86_tag <= cpu_tag;
        end
        if(_zz_863) begin
          ways_3_metas_87_tag <= cpu_tag;
        end
        if(_zz_864) begin
          ways_3_metas_88_tag <= cpu_tag;
        end
        if(_zz_865) begin
          ways_3_metas_89_tag <= cpu_tag;
        end
        if(_zz_866) begin
          ways_3_metas_90_tag <= cpu_tag;
        end
        if(_zz_867) begin
          ways_3_metas_91_tag <= cpu_tag;
        end
        if(_zz_868) begin
          ways_3_metas_92_tag <= cpu_tag;
        end
        if(_zz_869) begin
          ways_3_metas_93_tag <= cpu_tag;
        end
        if(_zz_870) begin
          ways_3_metas_94_tag <= cpu_tag;
        end
        if(_zz_871) begin
          ways_3_metas_95_tag <= cpu_tag;
        end
        if(_zz_872) begin
          ways_3_metas_96_tag <= cpu_tag;
        end
        if(_zz_873) begin
          ways_3_metas_97_tag <= cpu_tag;
        end
        if(_zz_874) begin
          ways_3_metas_98_tag <= cpu_tag;
        end
        if(_zz_875) begin
          ways_3_metas_99_tag <= cpu_tag;
        end
        if(_zz_876) begin
          ways_3_metas_100_tag <= cpu_tag;
        end
        if(_zz_877) begin
          ways_3_metas_101_tag <= cpu_tag;
        end
        if(_zz_878) begin
          ways_3_metas_102_tag <= cpu_tag;
        end
        if(_zz_879) begin
          ways_3_metas_103_tag <= cpu_tag;
        end
        if(_zz_880) begin
          ways_3_metas_104_tag <= cpu_tag;
        end
        if(_zz_881) begin
          ways_3_metas_105_tag <= cpu_tag;
        end
        if(_zz_882) begin
          ways_3_metas_106_tag <= cpu_tag;
        end
        if(_zz_883) begin
          ways_3_metas_107_tag <= cpu_tag;
        end
        if(_zz_884) begin
          ways_3_metas_108_tag <= cpu_tag;
        end
        if(_zz_885) begin
          ways_3_metas_109_tag <= cpu_tag;
        end
        if(_zz_886) begin
          ways_3_metas_110_tag <= cpu_tag;
        end
        if(_zz_887) begin
          ways_3_metas_111_tag <= cpu_tag;
        end
        if(_zz_888) begin
          ways_3_metas_112_tag <= cpu_tag;
        end
        if(_zz_889) begin
          ways_3_metas_113_tag <= cpu_tag;
        end
        if(_zz_890) begin
          ways_3_metas_114_tag <= cpu_tag;
        end
        if(_zz_891) begin
          ways_3_metas_115_tag <= cpu_tag;
        end
        if(_zz_892) begin
          ways_3_metas_116_tag <= cpu_tag;
        end
        if(_zz_893) begin
          ways_3_metas_117_tag <= cpu_tag;
        end
        if(_zz_894) begin
          ways_3_metas_118_tag <= cpu_tag;
        end
        if(_zz_895) begin
          ways_3_metas_119_tag <= cpu_tag;
        end
        if(_zz_896) begin
          ways_3_metas_120_tag <= cpu_tag;
        end
        if(_zz_897) begin
          ways_3_metas_121_tag <= cpu_tag;
        end
        if(_zz_898) begin
          ways_3_metas_122_tag <= cpu_tag;
        end
        if(_zz_899) begin
          ways_3_metas_123_tag <= cpu_tag;
        end
        if(_zz_900) begin
          ways_3_metas_124_tag <= cpu_tag;
        end
        if(_zz_901) begin
          ways_3_metas_125_tag <= cpu_tag;
        end
        if(_zz_902) begin
          ways_3_metas_126_tag <= cpu_tag;
        end
        if(_zz_903) begin
          ways_3_metas_127_tag <= cpu_tag;
        end
      end
      if(when_DCache_l237_3) begin
        cpu_cmd_ready_1 <= 1'b0;
      end else begin
        if(when_DCache_l240_3) begin
          cpu_cmd_ready_1 <= 1'b1;
        end
      end
    end
  end

  always @(posedge clk) begin
    if(is_miss) begin
      evict_id_miss <= evict_id;
    end
    next_level_rdone <= (next_level_rvalid && (next_level_data_cnt_value == 3'b111));
    next_level_wdone <= ((next_level_rsp_valid && (! next_level_rsp_payload_rvalid)) && (next_level_rsp_payload_bresp == 2'b00));
  end


endmodule

module SramBanks (
  input               sram_0_ports_cmd_valid,
  input      [6:0]    sram_0_ports_cmd_payload_addr,
  input      [15:0]   sram_0_ports_cmd_payload_wen,
  input      [511:0]  sram_0_ports_cmd_payload_wdata,
  input      [63:0]   sram_0_ports_cmd_payload_wstrb,
  output              sram_0_ports_rsp_valid,
  output reg [511:0]  sram_0_ports_rsp_payload_data,
  input               sram_1_ports_cmd_valid,
  input      [6:0]    sram_1_ports_cmd_payload_addr,
  input      [15:0]   sram_1_ports_cmd_payload_wen,
  input      [511:0]  sram_1_ports_cmd_payload_wdata,
  input      [63:0]   sram_1_ports_cmd_payload_wstrb,
  output              sram_1_ports_rsp_valid,
  output reg [511:0]  sram_1_ports_rsp_payload_data,
  input               sram_2_ports_cmd_valid,
  input      [6:0]    sram_2_ports_cmd_payload_addr,
  input      [15:0]   sram_2_ports_cmd_payload_wen,
  input      [511:0]  sram_2_ports_cmd_payload_wdata,
  input      [63:0]   sram_2_ports_cmd_payload_wstrb,
  output              sram_2_ports_rsp_valid,
  output reg [511:0]  sram_2_ports_rsp_payload_data,
  input               sram_3_ports_cmd_valid,
  input      [6:0]    sram_3_ports_cmd_payload_addr,
  input      [15:0]   sram_3_ports_cmd_payload_wen,
  input      [511:0]  sram_3_ports_cmd_payload_wdata,
  input      [63:0]   sram_3_ports_cmd_payload_wstrb,
  output              sram_3_ports_rsp_valid,
  output reg [511:0]  sram_3_ports_rsp_payload_data,
  input               clk,
  input               reset
);

  reg        [31:0]   _zz_sram_0_banks_0_bank_port1;
  reg        [31:0]   _zz_sram_0_banks_1_bank_port1;
  reg        [31:0]   _zz_sram_0_banks_2_bank_port1;
  reg        [31:0]   _zz_sram_0_banks_3_bank_port1;
  reg        [31:0]   _zz_sram_0_banks_4_bank_port1;
  reg        [31:0]   _zz_sram_0_banks_5_bank_port1;
  reg        [31:0]   _zz_sram_0_banks_6_bank_port1;
  reg        [31:0]   _zz_sram_0_banks_7_bank_port1;
  reg        [31:0]   _zz_sram_0_banks_8_bank_port1;
  reg        [31:0]   _zz_sram_0_banks_9_bank_port1;
  reg        [31:0]   _zz_sram_0_banks_10_bank_port1;
  reg        [31:0]   _zz_sram_0_banks_11_bank_port1;
  reg        [31:0]   _zz_sram_0_banks_12_bank_port1;
  reg        [31:0]   _zz_sram_0_banks_13_bank_port1;
  reg        [31:0]   _zz_sram_0_banks_14_bank_port1;
  reg        [31:0]   _zz_sram_0_banks_15_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_0_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_1_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_2_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_3_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_4_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_5_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_6_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_7_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_8_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_9_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_10_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_11_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_12_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_13_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_14_bank_port1;
  reg        [31:0]   _zz_sram_1_banks_15_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_0_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_1_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_2_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_3_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_4_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_5_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_6_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_7_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_8_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_9_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_10_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_11_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_12_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_13_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_14_bank_port1;
  reg        [31:0]   _zz_sram_2_banks_15_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_0_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_1_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_2_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_3_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_4_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_5_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_6_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_7_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_8_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_9_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_10_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_11_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_12_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_13_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_14_bank_port1;
  reg        [31:0]   _zz_sram_3_banks_15_bank_port1;
  wire       [31:0]   _zz_sram_0_banks_0_bank_port;
  wire       [3:0]    _zz_sram_0_banks_0_bank_port_1;
  wire                _zz_sram_0_banks_0_bank_port_2;
  wire       [31:0]   _zz_sram_0_banks_1_bank_port;
  wire       [3:0]    _zz_sram_0_banks_1_bank_port_1;
  wire                _zz_sram_0_banks_1_bank_port_2;
  wire       [31:0]   _zz_sram_0_banks_2_bank_port;
  wire       [3:0]    _zz_sram_0_banks_2_bank_port_1;
  wire                _zz_sram_0_banks_2_bank_port_2;
  wire       [31:0]   _zz_sram_0_banks_3_bank_port;
  wire       [3:0]    _zz_sram_0_banks_3_bank_port_1;
  wire                _zz_sram_0_banks_3_bank_port_2;
  wire       [31:0]   _zz_sram_0_banks_4_bank_port;
  wire       [3:0]    _zz_sram_0_banks_4_bank_port_1;
  wire                _zz_sram_0_banks_4_bank_port_2;
  wire       [31:0]   _zz_sram_0_banks_5_bank_port;
  wire       [3:0]    _zz_sram_0_banks_5_bank_port_1;
  wire                _zz_sram_0_banks_5_bank_port_2;
  wire       [31:0]   _zz_sram_0_banks_6_bank_port;
  wire       [3:0]    _zz_sram_0_banks_6_bank_port_1;
  wire                _zz_sram_0_banks_6_bank_port_2;
  wire       [31:0]   _zz_sram_0_banks_7_bank_port;
  wire       [3:0]    _zz_sram_0_banks_7_bank_port_1;
  wire                _zz_sram_0_banks_7_bank_port_2;
  wire       [31:0]   _zz_sram_0_banks_8_bank_port;
  wire       [3:0]    _zz_sram_0_banks_8_bank_port_1;
  wire                _zz_sram_0_banks_8_bank_port_2;
  wire       [31:0]   _zz_sram_0_banks_9_bank_port;
  wire       [3:0]    _zz_sram_0_banks_9_bank_port_1;
  wire                _zz_sram_0_banks_9_bank_port_2;
  wire       [31:0]   _zz_sram_0_banks_10_bank_port;
  wire       [3:0]    _zz_sram_0_banks_10_bank_port_1;
  wire                _zz_sram_0_banks_10_bank_port_2;
  wire       [31:0]   _zz_sram_0_banks_11_bank_port;
  wire       [3:0]    _zz_sram_0_banks_11_bank_port_1;
  wire                _zz_sram_0_banks_11_bank_port_2;
  wire       [31:0]   _zz_sram_0_banks_12_bank_port;
  wire       [3:0]    _zz_sram_0_banks_12_bank_port_1;
  wire                _zz_sram_0_banks_12_bank_port_2;
  wire       [31:0]   _zz_sram_0_banks_13_bank_port;
  wire       [3:0]    _zz_sram_0_banks_13_bank_port_1;
  wire                _zz_sram_0_banks_13_bank_port_2;
  wire       [31:0]   _zz_sram_0_banks_14_bank_port;
  wire       [3:0]    _zz_sram_0_banks_14_bank_port_1;
  wire                _zz_sram_0_banks_14_bank_port_2;
  wire       [31:0]   _zz_sram_0_banks_15_bank_port;
  wire       [3:0]    _zz_sram_0_banks_15_bank_port_1;
  wire                _zz_sram_0_banks_15_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_0_bank_port;
  wire       [3:0]    _zz_sram_1_banks_0_bank_port_1;
  wire                _zz_sram_1_banks_0_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_1_bank_port;
  wire       [3:0]    _zz_sram_1_banks_1_bank_port_1;
  wire                _zz_sram_1_banks_1_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_2_bank_port;
  wire       [3:0]    _zz_sram_1_banks_2_bank_port_1;
  wire                _zz_sram_1_banks_2_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_3_bank_port;
  wire       [3:0]    _zz_sram_1_banks_3_bank_port_1;
  wire                _zz_sram_1_banks_3_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_4_bank_port;
  wire       [3:0]    _zz_sram_1_banks_4_bank_port_1;
  wire                _zz_sram_1_banks_4_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_5_bank_port;
  wire       [3:0]    _zz_sram_1_banks_5_bank_port_1;
  wire                _zz_sram_1_banks_5_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_6_bank_port;
  wire       [3:0]    _zz_sram_1_banks_6_bank_port_1;
  wire                _zz_sram_1_banks_6_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_7_bank_port;
  wire       [3:0]    _zz_sram_1_banks_7_bank_port_1;
  wire                _zz_sram_1_banks_7_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_8_bank_port;
  wire       [3:0]    _zz_sram_1_banks_8_bank_port_1;
  wire                _zz_sram_1_banks_8_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_9_bank_port;
  wire       [3:0]    _zz_sram_1_banks_9_bank_port_1;
  wire                _zz_sram_1_banks_9_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_10_bank_port;
  wire       [3:0]    _zz_sram_1_banks_10_bank_port_1;
  wire                _zz_sram_1_banks_10_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_11_bank_port;
  wire       [3:0]    _zz_sram_1_banks_11_bank_port_1;
  wire                _zz_sram_1_banks_11_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_12_bank_port;
  wire       [3:0]    _zz_sram_1_banks_12_bank_port_1;
  wire                _zz_sram_1_banks_12_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_13_bank_port;
  wire       [3:0]    _zz_sram_1_banks_13_bank_port_1;
  wire                _zz_sram_1_banks_13_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_14_bank_port;
  wire       [3:0]    _zz_sram_1_banks_14_bank_port_1;
  wire                _zz_sram_1_banks_14_bank_port_2;
  wire       [31:0]   _zz_sram_1_banks_15_bank_port;
  wire       [3:0]    _zz_sram_1_banks_15_bank_port_1;
  wire                _zz_sram_1_banks_15_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_0_bank_port;
  wire       [3:0]    _zz_sram_2_banks_0_bank_port_1;
  wire                _zz_sram_2_banks_0_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_1_bank_port;
  wire       [3:0]    _zz_sram_2_banks_1_bank_port_1;
  wire                _zz_sram_2_banks_1_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_2_bank_port;
  wire       [3:0]    _zz_sram_2_banks_2_bank_port_1;
  wire                _zz_sram_2_banks_2_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_3_bank_port;
  wire       [3:0]    _zz_sram_2_banks_3_bank_port_1;
  wire                _zz_sram_2_banks_3_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_4_bank_port;
  wire       [3:0]    _zz_sram_2_banks_4_bank_port_1;
  wire                _zz_sram_2_banks_4_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_5_bank_port;
  wire       [3:0]    _zz_sram_2_banks_5_bank_port_1;
  wire                _zz_sram_2_banks_5_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_6_bank_port;
  wire       [3:0]    _zz_sram_2_banks_6_bank_port_1;
  wire                _zz_sram_2_banks_6_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_7_bank_port;
  wire       [3:0]    _zz_sram_2_banks_7_bank_port_1;
  wire                _zz_sram_2_banks_7_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_8_bank_port;
  wire       [3:0]    _zz_sram_2_banks_8_bank_port_1;
  wire                _zz_sram_2_banks_8_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_9_bank_port;
  wire       [3:0]    _zz_sram_2_banks_9_bank_port_1;
  wire                _zz_sram_2_banks_9_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_10_bank_port;
  wire       [3:0]    _zz_sram_2_banks_10_bank_port_1;
  wire                _zz_sram_2_banks_10_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_11_bank_port;
  wire       [3:0]    _zz_sram_2_banks_11_bank_port_1;
  wire                _zz_sram_2_banks_11_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_12_bank_port;
  wire       [3:0]    _zz_sram_2_banks_12_bank_port_1;
  wire                _zz_sram_2_banks_12_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_13_bank_port;
  wire       [3:0]    _zz_sram_2_banks_13_bank_port_1;
  wire                _zz_sram_2_banks_13_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_14_bank_port;
  wire       [3:0]    _zz_sram_2_banks_14_bank_port_1;
  wire                _zz_sram_2_banks_14_bank_port_2;
  wire       [31:0]   _zz_sram_2_banks_15_bank_port;
  wire       [3:0]    _zz_sram_2_banks_15_bank_port_1;
  wire                _zz_sram_2_banks_15_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_0_bank_port;
  wire       [3:0]    _zz_sram_3_banks_0_bank_port_1;
  wire                _zz_sram_3_banks_0_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_1_bank_port;
  wire       [3:0]    _zz_sram_3_banks_1_bank_port_1;
  wire                _zz_sram_3_banks_1_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_2_bank_port;
  wire       [3:0]    _zz_sram_3_banks_2_bank_port_1;
  wire                _zz_sram_3_banks_2_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_3_bank_port;
  wire       [3:0]    _zz_sram_3_banks_3_bank_port_1;
  wire                _zz_sram_3_banks_3_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_4_bank_port;
  wire       [3:0]    _zz_sram_3_banks_4_bank_port_1;
  wire                _zz_sram_3_banks_4_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_5_bank_port;
  wire       [3:0]    _zz_sram_3_banks_5_bank_port_1;
  wire                _zz_sram_3_banks_5_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_6_bank_port;
  wire       [3:0]    _zz_sram_3_banks_6_bank_port_1;
  wire                _zz_sram_3_banks_6_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_7_bank_port;
  wire       [3:0]    _zz_sram_3_banks_7_bank_port_1;
  wire                _zz_sram_3_banks_7_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_8_bank_port;
  wire       [3:0]    _zz_sram_3_banks_8_bank_port_1;
  wire                _zz_sram_3_banks_8_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_9_bank_port;
  wire       [3:0]    _zz_sram_3_banks_9_bank_port_1;
  wire                _zz_sram_3_banks_9_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_10_bank_port;
  wire       [3:0]    _zz_sram_3_banks_10_bank_port_1;
  wire                _zz_sram_3_banks_10_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_11_bank_port;
  wire       [3:0]    _zz_sram_3_banks_11_bank_port_1;
  wire                _zz_sram_3_banks_11_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_12_bank_port;
  wire       [3:0]    _zz_sram_3_banks_12_bank_port_1;
  wire                _zz_sram_3_banks_12_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_13_bank_port;
  wire       [3:0]    _zz_sram_3_banks_13_bank_port_1;
  wire                _zz_sram_3_banks_13_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_14_bank_port;
  wire       [3:0]    _zz_sram_3_banks_14_bank_port_1;
  wire                _zz_sram_3_banks_14_bank_port_2;
  wire       [31:0]   _zz_sram_3_banks_15_bank_port;
  wire       [3:0]    _zz_sram_3_banks_15_bank_port_1;
  wire                _zz_sram_3_banks_15_bank_port_2;
  reg                 _zz_sram_0_ports_rsp_valid;
  wire                when_SramBanks_l66;
  reg                 _zz_sram_1_ports_rsp_valid;
  wire                when_SramBanks_l66_1;
  reg                 _zz_sram_2_ports_rsp_valid;
  wire                when_SramBanks_l66_2;
  reg                 _zz_sram_3_ports_rsp_valid;
  wire                when_SramBanks_l66_3;
  reg [7:0] sram_0_banks_0_bank_symbol0 [0:127];
  reg [7:0] sram_0_banks_0_bank_symbol1 [0:127];
  reg [7:0] sram_0_banks_0_bank_symbol2 [0:127];
  reg [7:0] sram_0_banks_0_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_0_banks_0_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_0_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_0_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_0_banksymbol_read_3;
  reg [7:0] sram_0_banks_1_bank_symbol0 [0:127];
  reg [7:0] sram_0_banks_1_bank_symbol1 [0:127];
  reg [7:0] sram_0_banks_1_bank_symbol2 [0:127];
  reg [7:0] sram_0_banks_1_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_0_banks_1_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_1_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_1_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_1_banksymbol_read_3;
  reg [7:0] sram_0_banks_2_bank_symbol0 [0:127];
  reg [7:0] sram_0_banks_2_bank_symbol1 [0:127];
  reg [7:0] sram_0_banks_2_bank_symbol2 [0:127];
  reg [7:0] sram_0_banks_2_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_0_banks_2_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_2_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_2_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_2_banksymbol_read_3;
  reg [7:0] sram_0_banks_3_bank_symbol0 [0:127];
  reg [7:0] sram_0_banks_3_bank_symbol1 [0:127];
  reg [7:0] sram_0_banks_3_bank_symbol2 [0:127];
  reg [7:0] sram_0_banks_3_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_0_banks_3_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_3_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_3_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_3_banksymbol_read_3;
  reg [7:0] sram_0_banks_4_bank_symbol0 [0:127];
  reg [7:0] sram_0_banks_4_bank_symbol1 [0:127];
  reg [7:0] sram_0_banks_4_bank_symbol2 [0:127];
  reg [7:0] sram_0_banks_4_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_0_banks_4_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_4_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_4_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_4_banksymbol_read_3;
  reg [7:0] sram_0_banks_5_bank_symbol0 [0:127];
  reg [7:0] sram_0_banks_5_bank_symbol1 [0:127];
  reg [7:0] sram_0_banks_5_bank_symbol2 [0:127];
  reg [7:0] sram_0_banks_5_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_0_banks_5_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_5_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_5_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_5_banksymbol_read_3;
  reg [7:0] sram_0_banks_6_bank_symbol0 [0:127];
  reg [7:0] sram_0_banks_6_bank_symbol1 [0:127];
  reg [7:0] sram_0_banks_6_bank_symbol2 [0:127];
  reg [7:0] sram_0_banks_6_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_0_banks_6_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_6_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_6_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_6_banksymbol_read_3;
  reg [7:0] sram_0_banks_7_bank_symbol0 [0:127];
  reg [7:0] sram_0_banks_7_bank_symbol1 [0:127];
  reg [7:0] sram_0_banks_7_bank_symbol2 [0:127];
  reg [7:0] sram_0_banks_7_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_0_banks_7_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_7_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_7_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_7_banksymbol_read_3;
  reg [7:0] sram_0_banks_8_bank_symbol0 [0:127];
  reg [7:0] sram_0_banks_8_bank_symbol1 [0:127];
  reg [7:0] sram_0_banks_8_bank_symbol2 [0:127];
  reg [7:0] sram_0_banks_8_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_0_banks_8_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_8_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_8_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_8_banksymbol_read_3;
  reg [7:0] sram_0_banks_9_bank_symbol0 [0:127];
  reg [7:0] sram_0_banks_9_bank_symbol1 [0:127];
  reg [7:0] sram_0_banks_9_bank_symbol2 [0:127];
  reg [7:0] sram_0_banks_9_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_0_banks_9_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_9_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_9_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_9_banksymbol_read_3;
  reg [7:0] sram_0_banks_10_bank_symbol0 [0:127];
  reg [7:0] sram_0_banks_10_bank_symbol1 [0:127];
  reg [7:0] sram_0_banks_10_bank_symbol2 [0:127];
  reg [7:0] sram_0_banks_10_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_0_banks_10_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_10_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_10_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_10_banksymbol_read_3;
  reg [7:0] sram_0_banks_11_bank_symbol0 [0:127];
  reg [7:0] sram_0_banks_11_bank_symbol1 [0:127];
  reg [7:0] sram_0_banks_11_bank_symbol2 [0:127];
  reg [7:0] sram_0_banks_11_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_0_banks_11_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_11_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_11_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_11_banksymbol_read_3;
  reg [7:0] sram_0_banks_12_bank_symbol0 [0:127];
  reg [7:0] sram_0_banks_12_bank_symbol1 [0:127];
  reg [7:0] sram_0_banks_12_bank_symbol2 [0:127];
  reg [7:0] sram_0_banks_12_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_0_banks_12_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_12_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_12_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_12_banksymbol_read_3;
  reg [7:0] sram_0_banks_13_bank_symbol0 [0:127];
  reg [7:0] sram_0_banks_13_bank_symbol1 [0:127];
  reg [7:0] sram_0_banks_13_bank_symbol2 [0:127];
  reg [7:0] sram_0_banks_13_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_0_banks_13_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_13_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_13_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_13_banksymbol_read_3;
  reg [7:0] sram_0_banks_14_bank_symbol0 [0:127];
  reg [7:0] sram_0_banks_14_bank_symbol1 [0:127];
  reg [7:0] sram_0_banks_14_bank_symbol2 [0:127];
  reg [7:0] sram_0_banks_14_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_0_banks_14_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_14_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_14_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_14_banksymbol_read_3;
  reg [7:0] sram_0_banks_15_bank_symbol0 [0:127];
  reg [7:0] sram_0_banks_15_bank_symbol1 [0:127];
  reg [7:0] sram_0_banks_15_bank_symbol2 [0:127];
  reg [7:0] sram_0_banks_15_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_0_banks_15_banksymbol_read;
  reg [7:0] _zz_sram_0_banks_15_banksymbol_read_1;
  reg [7:0] _zz_sram_0_banks_15_banksymbol_read_2;
  reg [7:0] _zz_sram_0_banks_15_banksymbol_read_3;
  reg [7:0] sram_1_banks_0_bank_symbol0 [0:127];
  reg [7:0] sram_1_banks_0_bank_symbol1 [0:127];
  reg [7:0] sram_1_banks_0_bank_symbol2 [0:127];
  reg [7:0] sram_1_banks_0_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_1_banks_0_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_0_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_0_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_0_banksymbol_read_3;
  reg [7:0] sram_1_banks_1_bank_symbol0 [0:127];
  reg [7:0] sram_1_banks_1_bank_symbol1 [0:127];
  reg [7:0] sram_1_banks_1_bank_symbol2 [0:127];
  reg [7:0] sram_1_banks_1_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_1_banks_1_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_1_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_1_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_1_banksymbol_read_3;
  reg [7:0] sram_1_banks_2_bank_symbol0 [0:127];
  reg [7:0] sram_1_banks_2_bank_symbol1 [0:127];
  reg [7:0] sram_1_banks_2_bank_symbol2 [0:127];
  reg [7:0] sram_1_banks_2_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_1_banks_2_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_2_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_2_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_2_banksymbol_read_3;
  reg [7:0] sram_1_banks_3_bank_symbol0 [0:127];
  reg [7:0] sram_1_banks_3_bank_symbol1 [0:127];
  reg [7:0] sram_1_banks_3_bank_symbol2 [0:127];
  reg [7:0] sram_1_banks_3_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_1_banks_3_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_3_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_3_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_3_banksymbol_read_3;
  reg [7:0] sram_1_banks_4_bank_symbol0 [0:127];
  reg [7:0] sram_1_banks_4_bank_symbol1 [0:127];
  reg [7:0] sram_1_banks_4_bank_symbol2 [0:127];
  reg [7:0] sram_1_banks_4_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_1_banks_4_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_4_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_4_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_4_banksymbol_read_3;
  reg [7:0] sram_1_banks_5_bank_symbol0 [0:127];
  reg [7:0] sram_1_banks_5_bank_symbol1 [0:127];
  reg [7:0] sram_1_banks_5_bank_symbol2 [0:127];
  reg [7:0] sram_1_banks_5_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_1_banks_5_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_5_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_5_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_5_banksymbol_read_3;
  reg [7:0] sram_1_banks_6_bank_symbol0 [0:127];
  reg [7:0] sram_1_banks_6_bank_symbol1 [0:127];
  reg [7:0] sram_1_banks_6_bank_symbol2 [0:127];
  reg [7:0] sram_1_banks_6_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_1_banks_6_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_6_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_6_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_6_banksymbol_read_3;
  reg [7:0] sram_1_banks_7_bank_symbol0 [0:127];
  reg [7:0] sram_1_banks_7_bank_symbol1 [0:127];
  reg [7:0] sram_1_banks_7_bank_symbol2 [0:127];
  reg [7:0] sram_1_banks_7_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_1_banks_7_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_7_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_7_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_7_banksymbol_read_3;
  reg [7:0] sram_1_banks_8_bank_symbol0 [0:127];
  reg [7:0] sram_1_banks_8_bank_symbol1 [0:127];
  reg [7:0] sram_1_banks_8_bank_symbol2 [0:127];
  reg [7:0] sram_1_banks_8_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_1_banks_8_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_8_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_8_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_8_banksymbol_read_3;
  reg [7:0] sram_1_banks_9_bank_symbol0 [0:127];
  reg [7:0] sram_1_banks_9_bank_symbol1 [0:127];
  reg [7:0] sram_1_banks_9_bank_symbol2 [0:127];
  reg [7:0] sram_1_banks_9_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_1_banks_9_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_9_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_9_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_9_banksymbol_read_3;
  reg [7:0] sram_1_banks_10_bank_symbol0 [0:127];
  reg [7:0] sram_1_banks_10_bank_symbol1 [0:127];
  reg [7:0] sram_1_banks_10_bank_symbol2 [0:127];
  reg [7:0] sram_1_banks_10_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_1_banks_10_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_10_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_10_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_10_banksymbol_read_3;
  reg [7:0] sram_1_banks_11_bank_symbol0 [0:127];
  reg [7:0] sram_1_banks_11_bank_symbol1 [0:127];
  reg [7:0] sram_1_banks_11_bank_symbol2 [0:127];
  reg [7:0] sram_1_banks_11_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_1_banks_11_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_11_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_11_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_11_banksymbol_read_3;
  reg [7:0] sram_1_banks_12_bank_symbol0 [0:127];
  reg [7:0] sram_1_banks_12_bank_symbol1 [0:127];
  reg [7:0] sram_1_banks_12_bank_symbol2 [0:127];
  reg [7:0] sram_1_banks_12_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_1_banks_12_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_12_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_12_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_12_banksymbol_read_3;
  reg [7:0] sram_1_banks_13_bank_symbol0 [0:127];
  reg [7:0] sram_1_banks_13_bank_symbol1 [0:127];
  reg [7:0] sram_1_banks_13_bank_symbol2 [0:127];
  reg [7:0] sram_1_banks_13_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_1_banks_13_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_13_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_13_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_13_banksymbol_read_3;
  reg [7:0] sram_1_banks_14_bank_symbol0 [0:127];
  reg [7:0] sram_1_banks_14_bank_symbol1 [0:127];
  reg [7:0] sram_1_banks_14_bank_symbol2 [0:127];
  reg [7:0] sram_1_banks_14_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_1_banks_14_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_14_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_14_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_14_banksymbol_read_3;
  reg [7:0] sram_1_banks_15_bank_symbol0 [0:127];
  reg [7:0] sram_1_banks_15_bank_symbol1 [0:127];
  reg [7:0] sram_1_banks_15_bank_symbol2 [0:127];
  reg [7:0] sram_1_banks_15_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_1_banks_15_banksymbol_read;
  reg [7:0] _zz_sram_1_banks_15_banksymbol_read_1;
  reg [7:0] _zz_sram_1_banks_15_banksymbol_read_2;
  reg [7:0] _zz_sram_1_banks_15_banksymbol_read_3;
  reg [7:0] sram_2_banks_0_bank_symbol0 [0:127];
  reg [7:0] sram_2_banks_0_bank_symbol1 [0:127];
  reg [7:0] sram_2_banks_0_bank_symbol2 [0:127];
  reg [7:0] sram_2_banks_0_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_2_banks_0_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_0_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_0_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_0_banksymbol_read_3;
  reg [7:0] sram_2_banks_1_bank_symbol0 [0:127];
  reg [7:0] sram_2_banks_1_bank_symbol1 [0:127];
  reg [7:0] sram_2_banks_1_bank_symbol2 [0:127];
  reg [7:0] sram_2_banks_1_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_2_banks_1_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_1_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_1_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_1_banksymbol_read_3;
  reg [7:0] sram_2_banks_2_bank_symbol0 [0:127];
  reg [7:0] sram_2_banks_2_bank_symbol1 [0:127];
  reg [7:0] sram_2_banks_2_bank_symbol2 [0:127];
  reg [7:0] sram_2_banks_2_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_2_banks_2_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_2_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_2_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_2_banksymbol_read_3;
  reg [7:0] sram_2_banks_3_bank_symbol0 [0:127];
  reg [7:0] sram_2_banks_3_bank_symbol1 [0:127];
  reg [7:0] sram_2_banks_3_bank_symbol2 [0:127];
  reg [7:0] sram_2_banks_3_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_2_banks_3_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_3_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_3_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_3_banksymbol_read_3;
  reg [7:0] sram_2_banks_4_bank_symbol0 [0:127];
  reg [7:0] sram_2_banks_4_bank_symbol1 [0:127];
  reg [7:0] sram_2_banks_4_bank_symbol2 [0:127];
  reg [7:0] sram_2_banks_4_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_2_banks_4_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_4_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_4_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_4_banksymbol_read_3;
  reg [7:0] sram_2_banks_5_bank_symbol0 [0:127];
  reg [7:0] sram_2_banks_5_bank_symbol1 [0:127];
  reg [7:0] sram_2_banks_5_bank_symbol2 [0:127];
  reg [7:0] sram_2_banks_5_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_2_banks_5_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_5_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_5_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_5_banksymbol_read_3;
  reg [7:0] sram_2_banks_6_bank_symbol0 [0:127];
  reg [7:0] sram_2_banks_6_bank_symbol1 [0:127];
  reg [7:0] sram_2_banks_6_bank_symbol2 [0:127];
  reg [7:0] sram_2_banks_6_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_2_banks_6_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_6_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_6_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_6_banksymbol_read_3;
  reg [7:0] sram_2_banks_7_bank_symbol0 [0:127];
  reg [7:0] sram_2_banks_7_bank_symbol1 [0:127];
  reg [7:0] sram_2_banks_7_bank_symbol2 [0:127];
  reg [7:0] sram_2_banks_7_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_2_banks_7_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_7_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_7_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_7_banksymbol_read_3;
  reg [7:0] sram_2_banks_8_bank_symbol0 [0:127];
  reg [7:0] sram_2_banks_8_bank_symbol1 [0:127];
  reg [7:0] sram_2_banks_8_bank_symbol2 [0:127];
  reg [7:0] sram_2_banks_8_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_2_banks_8_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_8_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_8_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_8_banksymbol_read_3;
  reg [7:0] sram_2_banks_9_bank_symbol0 [0:127];
  reg [7:0] sram_2_banks_9_bank_symbol1 [0:127];
  reg [7:0] sram_2_banks_9_bank_symbol2 [0:127];
  reg [7:0] sram_2_banks_9_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_2_banks_9_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_9_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_9_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_9_banksymbol_read_3;
  reg [7:0] sram_2_banks_10_bank_symbol0 [0:127];
  reg [7:0] sram_2_banks_10_bank_symbol1 [0:127];
  reg [7:0] sram_2_banks_10_bank_symbol2 [0:127];
  reg [7:0] sram_2_banks_10_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_2_banks_10_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_10_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_10_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_10_banksymbol_read_3;
  reg [7:0] sram_2_banks_11_bank_symbol0 [0:127];
  reg [7:0] sram_2_banks_11_bank_symbol1 [0:127];
  reg [7:0] sram_2_banks_11_bank_symbol2 [0:127];
  reg [7:0] sram_2_banks_11_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_2_banks_11_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_11_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_11_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_11_banksymbol_read_3;
  reg [7:0] sram_2_banks_12_bank_symbol0 [0:127];
  reg [7:0] sram_2_banks_12_bank_symbol1 [0:127];
  reg [7:0] sram_2_banks_12_bank_symbol2 [0:127];
  reg [7:0] sram_2_banks_12_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_2_banks_12_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_12_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_12_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_12_banksymbol_read_3;
  reg [7:0] sram_2_banks_13_bank_symbol0 [0:127];
  reg [7:0] sram_2_banks_13_bank_symbol1 [0:127];
  reg [7:0] sram_2_banks_13_bank_symbol2 [0:127];
  reg [7:0] sram_2_banks_13_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_2_banks_13_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_13_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_13_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_13_banksymbol_read_3;
  reg [7:0] sram_2_banks_14_bank_symbol0 [0:127];
  reg [7:0] sram_2_banks_14_bank_symbol1 [0:127];
  reg [7:0] sram_2_banks_14_bank_symbol2 [0:127];
  reg [7:0] sram_2_banks_14_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_2_banks_14_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_14_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_14_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_14_banksymbol_read_3;
  reg [7:0] sram_2_banks_15_bank_symbol0 [0:127];
  reg [7:0] sram_2_banks_15_bank_symbol1 [0:127];
  reg [7:0] sram_2_banks_15_bank_symbol2 [0:127];
  reg [7:0] sram_2_banks_15_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_2_banks_15_banksymbol_read;
  reg [7:0] _zz_sram_2_banks_15_banksymbol_read_1;
  reg [7:0] _zz_sram_2_banks_15_banksymbol_read_2;
  reg [7:0] _zz_sram_2_banks_15_banksymbol_read_3;
  reg [7:0] sram_3_banks_0_bank_symbol0 [0:127];
  reg [7:0] sram_3_banks_0_bank_symbol1 [0:127];
  reg [7:0] sram_3_banks_0_bank_symbol2 [0:127];
  reg [7:0] sram_3_banks_0_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_3_banks_0_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_0_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_0_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_0_banksymbol_read_3;
  reg [7:0] sram_3_banks_1_bank_symbol0 [0:127];
  reg [7:0] sram_3_banks_1_bank_symbol1 [0:127];
  reg [7:0] sram_3_banks_1_bank_symbol2 [0:127];
  reg [7:0] sram_3_banks_1_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_3_banks_1_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_1_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_1_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_1_banksymbol_read_3;
  reg [7:0] sram_3_banks_2_bank_symbol0 [0:127];
  reg [7:0] sram_3_banks_2_bank_symbol1 [0:127];
  reg [7:0] sram_3_banks_2_bank_symbol2 [0:127];
  reg [7:0] sram_3_banks_2_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_3_banks_2_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_2_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_2_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_2_banksymbol_read_3;
  reg [7:0] sram_3_banks_3_bank_symbol0 [0:127];
  reg [7:0] sram_3_banks_3_bank_symbol1 [0:127];
  reg [7:0] sram_3_banks_3_bank_symbol2 [0:127];
  reg [7:0] sram_3_banks_3_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_3_banks_3_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_3_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_3_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_3_banksymbol_read_3;
  reg [7:0] sram_3_banks_4_bank_symbol0 [0:127];
  reg [7:0] sram_3_banks_4_bank_symbol1 [0:127];
  reg [7:0] sram_3_banks_4_bank_symbol2 [0:127];
  reg [7:0] sram_3_banks_4_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_3_banks_4_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_4_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_4_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_4_banksymbol_read_3;
  reg [7:0] sram_3_banks_5_bank_symbol0 [0:127];
  reg [7:0] sram_3_banks_5_bank_symbol1 [0:127];
  reg [7:0] sram_3_banks_5_bank_symbol2 [0:127];
  reg [7:0] sram_3_banks_5_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_3_banks_5_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_5_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_5_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_5_banksymbol_read_3;
  reg [7:0] sram_3_banks_6_bank_symbol0 [0:127];
  reg [7:0] sram_3_banks_6_bank_symbol1 [0:127];
  reg [7:0] sram_3_banks_6_bank_symbol2 [0:127];
  reg [7:0] sram_3_banks_6_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_3_banks_6_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_6_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_6_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_6_banksymbol_read_3;
  reg [7:0] sram_3_banks_7_bank_symbol0 [0:127];
  reg [7:0] sram_3_banks_7_bank_symbol1 [0:127];
  reg [7:0] sram_3_banks_7_bank_symbol2 [0:127];
  reg [7:0] sram_3_banks_7_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_3_banks_7_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_7_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_7_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_7_banksymbol_read_3;
  reg [7:0] sram_3_banks_8_bank_symbol0 [0:127];
  reg [7:0] sram_3_banks_8_bank_symbol1 [0:127];
  reg [7:0] sram_3_banks_8_bank_symbol2 [0:127];
  reg [7:0] sram_3_banks_8_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_3_banks_8_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_8_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_8_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_8_banksymbol_read_3;
  reg [7:0] sram_3_banks_9_bank_symbol0 [0:127];
  reg [7:0] sram_3_banks_9_bank_symbol1 [0:127];
  reg [7:0] sram_3_banks_9_bank_symbol2 [0:127];
  reg [7:0] sram_3_banks_9_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_3_banks_9_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_9_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_9_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_9_banksymbol_read_3;
  reg [7:0] sram_3_banks_10_bank_symbol0 [0:127];
  reg [7:0] sram_3_banks_10_bank_symbol1 [0:127];
  reg [7:0] sram_3_banks_10_bank_symbol2 [0:127];
  reg [7:0] sram_3_banks_10_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_3_banks_10_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_10_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_10_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_10_banksymbol_read_3;
  reg [7:0] sram_3_banks_11_bank_symbol0 [0:127];
  reg [7:0] sram_3_banks_11_bank_symbol1 [0:127];
  reg [7:0] sram_3_banks_11_bank_symbol2 [0:127];
  reg [7:0] sram_3_banks_11_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_3_banks_11_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_11_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_11_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_11_banksymbol_read_3;
  reg [7:0] sram_3_banks_12_bank_symbol0 [0:127];
  reg [7:0] sram_3_banks_12_bank_symbol1 [0:127];
  reg [7:0] sram_3_banks_12_bank_symbol2 [0:127];
  reg [7:0] sram_3_banks_12_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_3_banks_12_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_12_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_12_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_12_banksymbol_read_3;
  reg [7:0] sram_3_banks_13_bank_symbol0 [0:127];
  reg [7:0] sram_3_banks_13_bank_symbol1 [0:127];
  reg [7:0] sram_3_banks_13_bank_symbol2 [0:127];
  reg [7:0] sram_3_banks_13_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_3_banks_13_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_13_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_13_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_13_banksymbol_read_3;
  reg [7:0] sram_3_banks_14_bank_symbol0 [0:127];
  reg [7:0] sram_3_banks_14_bank_symbol1 [0:127];
  reg [7:0] sram_3_banks_14_bank_symbol2 [0:127];
  reg [7:0] sram_3_banks_14_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_3_banks_14_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_14_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_14_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_14_banksymbol_read_3;
  reg [7:0] sram_3_banks_15_bank_symbol0 [0:127];
  reg [7:0] sram_3_banks_15_bank_symbol1 [0:127];
  reg [7:0] sram_3_banks_15_bank_symbol2 [0:127];
  reg [7:0] sram_3_banks_15_bank_symbol3 [0:127];
  reg [7:0] _zz_sram_3_banks_15_banksymbol_read;
  reg [7:0] _zz_sram_3_banks_15_banksymbol_read_1;
  reg [7:0] _zz_sram_3_banks_15_banksymbol_read_2;
  reg [7:0] _zz_sram_3_banks_15_banksymbol_read_3;

  assign _zz_sram_0_banks_0_bank_port = sram_0_ports_cmd_payload_wdata[31 : 0];
  assign _zz_sram_0_banks_0_bank_port_1 = sram_0_ports_cmd_payload_wstrb[3 : 0];
  assign _zz_sram_0_banks_0_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[0]);
  assign _zz_sram_0_banks_1_bank_port = sram_0_ports_cmd_payload_wdata[63 : 32];
  assign _zz_sram_0_banks_1_bank_port_1 = sram_0_ports_cmd_payload_wstrb[7 : 4];
  assign _zz_sram_0_banks_1_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[1]);
  assign _zz_sram_0_banks_2_bank_port = sram_0_ports_cmd_payload_wdata[95 : 64];
  assign _zz_sram_0_banks_2_bank_port_1 = sram_0_ports_cmd_payload_wstrb[11 : 8];
  assign _zz_sram_0_banks_2_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[2]);
  assign _zz_sram_0_banks_3_bank_port = sram_0_ports_cmd_payload_wdata[127 : 96];
  assign _zz_sram_0_banks_3_bank_port_1 = sram_0_ports_cmd_payload_wstrb[15 : 12];
  assign _zz_sram_0_banks_3_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[3]);
  assign _zz_sram_0_banks_4_bank_port = sram_0_ports_cmd_payload_wdata[159 : 128];
  assign _zz_sram_0_banks_4_bank_port_1 = sram_0_ports_cmd_payload_wstrb[19 : 16];
  assign _zz_sram_0_banks_4_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[4]);
  assign _zz_sram_0_banks_5_bank_port = sram_0_ports_cmd_payload_wdata[191 : 160];
  assign _zz_sram_0_banks_5_bank_port_1 = sram_0_ports_cmd_payload_wstrb[23 : 20];
  assign _zz_sram_0_banks_5_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[5]);
  assign _zz_sram_0_banks_6_bank_port = sram_0_ports_cmd_payload_wdata[223 : 192];
  assign _zz_sram_0_banks_6_bank_port_1 = sram_0_ports_cmd_payload_wstrb[27 : 24];
  assign _zz_sram_0_banks_6_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[6]);
  assign _zz_sram_0_banks_7_bank_port = sram_0_ports_cmd_payload_wdata[255 : 224];
  assign _zz_sram_0_banks_7_bank_port_1 = sram_0_ports_cmd_payload_wstrb[31 : 28];
  assign _zz_sram_0_banks_7_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[7]);
  assign _zz_sram_0_banks_8_bank_port = sram_0_ports_cmd_payload_wdata[287 : 256];
  assign _zz_sram_0_banks_8_bank_port_1 = sram_0_ports_cmd_payload_wstrb[35 : 32];
  assign _zz_sram_0_banks_8_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[8]);
  assign _zz_sram_0_banks_9_bank_port = sram_0_ports_cmd_payload_wdata[319 : 288];
  assign _zz_sram_0_banks_9_bank_port_1 = sram_0_ports_cmd_payload_wstrb[39 : 36];
  assign _zz_sram_0_banks_9_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[9]);
  assign _zz_sram_0_banks_10_bank_port = sram_0_ports_cmd_payload_wdata[351 : 320];
  assign _zz_sram_0_banks_10_bank_port_1 = sram_0_ports_cmd_payload_wstrb[43 : 40];
  assign _zz_sram_0_banks_10_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[10]);
  assign _zz_sram_0_banks_11_bank_port = sram_0_ports_cmd_payload_wdata[383 : 352];
  assign _zz_sram_0_banks_11_bank_port_1 = sram_0_ports_cmd_payload_wstrb[47 : 44];
  assign _zz_sram_0_banks_11_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[11]);
  assign _zz_sram_0_banks_12_bank_port = sram_0_ports_cmd_payload_wdata[415 : 384];
  assign _zz_sram_0_banks_12_bank_port_1 = sram_0_ports_cmd_payload_wstrb[51 : 48];
  assign _zz_sram_0_banks_12_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[12]);
  assign _zz_sram_0_banks_13_bank_port = sram_0_ports_cmd_payload_wdata[447 : 416];
  assign _zz_sram_0_banks_13_bank_port_1 = sram_0_ports_cmd_payload_wstrb[55 : 52];
  assign _zz_sram_0_banks_13_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[13]);
  assign _zz_sram_0_banks_14_bank_port = sram_0_ports_cmd_payload_wdata[479 : 448];
  assign _zz_sram_0_banks_14_bank_port_1 = sram_0_ports_cmd_payload_wstrb[59 : 56];
  assign _zz_sram_0_banks_14_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[14]);
  assign _zz_sram_0_banks_15_bank_port = sram_0_ports_cmd_payload_wdata[511 : 480];
  assign _zz_sram_0_banks_15_bank_port_1 = sram_0_ports_cmd_payload_wstrb[63 : 60];
  assign _zz_sram_0_banks_15_bank_port_2 = (sram_0_ports_cmd_valid && sram_0_ports_cmd_payload_wen[15]);
  assign _zz_sram_1_banks_0_bank_port = sram_1_ports_cmd_payload_wdata[31 : 0];
  assign _zz_sram_1_banks_0_bank_port_1 = sram_1_ports_cmd_payload_wstrb[3 : 0];
  assign _zz_sram_1_banks_0_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[0]);
  assign _zz_sram_1_banks_1_bank_port = sram_1_ports_cmd_payload_wdata[63 : 32];
  assign _zz_sram_1_banks_1_bank_port_1 = sram_1_ports_cmd_payload_wstrb[7 : 4];
  assign _zz_sram_1_banks_1_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[1]);
  assign _zz_sram_1_banks_2_bank_port = sram_1_ports_cmd_payload_wdata[95 : 64];
  assign _zz_sram_1_banks_2_bank_port_1 = sram_1_ports_cmd_payload_wstrb[11 : 8];
  assign _zz_sram_1_banks_2_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[2]);
  assign _zz_sram_1_banks_3_bank_port = sram_1_ports_cmd_payload_wdata[127 : 96];
  assign _zz_sram_1_banks_3_bank_port_1 = sram_1_ports_cmd_payload_wstrb[15 : 12];
  assign _zz_sram_1_banks_3_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[3]);
  assign _zz_sram_1_banks_4_bank_port = sram_1_ports_cmd_payload_wdata[159 : 128];
  assign _zz_sram_1_banks_4_bank_port_1 = sram_1_ports_cmd_payload_wstrb[19 : 16];
  assign _zz_sram_1_banks_4_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[4]);
  assign _zz_sram_1_banks_5_bank_port = sram_1_ports_cmd_payload_wdata[191 : 160];
  assign _zz_sram_1_banks_5_bank_port_1 = sram_1_ports_cmd_payload_wstrb[23 : 20];
  assign _zz_sram_1_banks_5_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[5]);
  assign _zz_sram_1_banks_6_bank_port = sram_1_ports_cmd_payload_wdata[223 : 192];
  assign _zz_sram_1_banks_6_bank_port_1 = sram_1_ports_cmd_payload_wstrb[27 : 24];
  assign _zz_sram_1_banks_6_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[6]);
  assign _zz_sram_1_banks_7_bank_port = sram_1_ports_cmd_payload_wdata[255 : 224];
  assign _zz_sram_1_banks_7_bank_port_1 = sram_1_ports_cmd_payload_wstrb[31 : 28];
  assign _zz_sram_1_banks_7_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[7]);
  assign _zz_sram_1_banks_8_bank_port = sram_1_ports_cmd_payload_wdata[287 : 256];
  assign _zz_sram_1_banks_8_bank_port_1 = sram_1_ports_cmd_payload_wstrb[35 : 32];
  assign _zz_sram_1_banks_8_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[8]);
  assign _zz_sram_1_banks_9_bank_port = sram_1_ports_cmd_payload_wdata[319 : 288];
  assign _zz_sram_1_banks_9_bank_port_1 = sram_1_ports_cmd_payload_wstrb[39 : 36];
  assign _zz_sram_1_banks_9_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[9]);
  assign _zz_sram_1_banks_10_bank_port = sram_1_ports_cmd_payload_wdata[351 : 320];
  assign _zz_sram_1_banks_10_bank_port_1 = sram_1_ports_cmd_payload_wstrb[43 : 40];
  assign _zz_sram_1_banks_10_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[10]);
  assign _zz_sram_1_banks_11_bank_port = sram_1_ports_cmd_payload_wdata[383 : 352];
  assign _zz_sram_1_banks_11_bank_port_1 = sram_1_ports_cmd_payload_wstrb[47 : 44];
  assign _zz_sram_1_banks_11_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[11]);
  assign _zz_sram_1_banks_12_bank_port = sram_1_ports_cmd_payload_wdata[415 : 384];
  assign _zz_sram_1_banks_12_bank_port_1 = sram_1_ports_cmd_payload_wstrb[51 : 48];
  assign _zz_sram_1_banks_12_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[12]);
  assign _zz_sram_1_banks_13_bank_port = sram_1_ports_cmd_payload_wdata[447 : 416];
  assign _zz_sram_1_banks_13_bank_port_1 = sram_1_ports_cmd_payload_wstrb[55 : 52];
  assign _zz_sram_1_banks_13_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[13]);
  assign _zz_sram_1_banks_14_bank_port = sram_1_ports_cmd_payload_wdata[479 : 448];
  assign _zz_sram_1_banks_14_bank_port_1 = sram_1_ports_cmd_payload_wstrb[59 : 56];
  assign _zz_sram_1_banks_14_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[14]);
  assign _zz_sram_1_banks_15_bank_port = sram_1_ports_cmd_payload_wdata[511 : 480];
  assign _zz_sram_1_banks_15_bank_port_1 = sram_1_ports_cmd_payload_wstrb[63 : 60];
  assign _zz_sram_1_banks_15_bank_port_2 = (sram_1_ports_cmd_valid && sram_1_ports_cmd_payload_wen[15]);
  assign _zz_sram_2_banks_0_bank_port = sram_2_ports_cmd_payload_wdata[31 : 0];
  assign _zz_sram_2_banks_0_bank_port_1 = sram_2_ports_cmd_payload_wstrb[3 : 0];
  assign _zz_sram_2_banks_0_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[0]);
  assign _zz_sram_2_banks_1_bank_port = sram_2_ports_cmd_payload_wdata[63 : 32];
  assign _zz_sram_2_banks_1_bank_port_1 = sram_2_ports_cmd_payload_wstrb[7 : 4];
  assign _zz_sram_2_banks_1_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[1]);
  assign _zz_sram_2_banks_2_bank_port = sram_2_ports_cmd_payload_wdata[95 : 64];
  assign _zz_sram_2_banks_2_bank_port_1 = sram_2_ports_cmd_payload_wstrb[11 : 8];
  assign _zz_sram_2_banks_2_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[2]);
  assign _zz_sram_2_banks_3_bank_port = sram_2_ports_cmd_payload_wdata[127 : 96];
  assign _zz_sram_2_banks_3_bank_port_1 = sram_2_ports_cmd_payload_wstrb[15 : 12];
  assign _zz_sram_2_banks_3_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[3]);
  assign _zz_sram_2_banks_4_bank_port = sram_2_ports_cmd_payload_wdata[159 : 128];
  assign _zz_sram_2_banks_4_bank_port_1 = sram_2_ports_cmd_payload_wstrb[19 : 16];
  assign _zz_sram_2_banks_4_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[4]);
  assign _zz_sram_2_banks_5_bank_port = sram_2_ports_cmd_payload_wdata[191 : 160];
  assign _zz_sram_2_banks_5_bank_port_1 = sram_2_ports_cmd_payload_wstrb[23 : 20];
  assign _zz_sram_2_banks_5_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[5]);
  assign _zz_sram_2_banks_6_bank_port = sram_2_ports_cmd_payload_wdata[223 : 192];
  assign _zz_sram_2_banks_6_bank_port_1 = sram_2_ports_cmd_payload_wstrb[27 : 24];
  assign _zz_sram_2_banks_6_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[6]);
  assign _zz_sram_2_banks_7_bank_port = sram_2_ports_cmd_payload_wdata[255 : 224];
  assign _zz_sram_2_banks_7_bank_port_1 = sram_2_ports_cmd_payload_wstrb[31 : 28];
  assign _zz_sram_2_banks_7_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[7]);
  assign _zz_sram_2_banks_8_bank_port = sram_2_ports_cmd_payload_wdata[287 : 256];
  assign _zz_sram_2_banks_8_bank_port_1 = sram_2_ports_cmd_payload_wstrb[35 : 32];
  assign _zz_sram_2_banks_8_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[8]);
  assign _zz_sram_2_banks_9_bank_port = sram_2_ports_cmd_payload_wdata[319 : 288];
  assign _zz_sram_2_banks_9_bank_port_1 = sram_2_ports_cmd_payload_wstrb[39 : 36];
  assign _zz_sram_2_banks_9_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[9]);
  assign _zz_sram_2_banks_10_bank_port = sram_2_ports_cmd_payload_wdata[351 : 320];
  assign _zz_sram_2_banks_10_bank_port_1 = sram_2_ports_cmd_payload_wstrb[43 : 40];
  assign _zz_sram_2_banks_10_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[10]);
  assign _zz_sram_2_banks_11_bank_port = sram_2_ports_cmd_payload_wdata[383 : 352];
  assign _zz_sram_2_banks_11_bank_port_1 = sram_2_ports_cmd_payload_wstrb[47 : 44];
  assign _zz_sram_2_banks_11_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[11]);
  assign _zz_sram_2_banks_12_bank_port = sram_2_ports_cmd_payload_wdata[415 : 384];
  assign _zz_sram_2_banks_12_bank_port_1 = sram_2_ports_cmd_payload_wstrb[51 : 48];
  assign _zz_sram_2_banks_12_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[12]);
  assign _zz_sram_2_banks_13_bank_port = sram_2_ports_cmd_payload_wdata[447 : 416];
  assign _zz_sram_2_banks_13_bank_port_1 = sram_2_ports_cmd_payload_wstrb[55 : 52];
  assign _zz_sram_2_banks_13_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[13]);
  assign _zz_sram_2_banks_14_bank_port = sram_2_ports_cmd_payload_wdata[479 : 448];
  assign _zz_sram_2_banks_14_bank_port_1 = sram_2_ports_cmd_payload_wstrb[59 : 56];
  assign _zz_sram_2_banks_14_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[14]);
  assign _zz_sram_2_banks_15_bank_port = sram_2_ports_cmd_payload_wdata[511 : 480];
  assign _zz_sram_2_banks_15_bank_port_1 = sram_2_ports_cmd_payload_wstrb[63 : 60];
  assign _zz_sram_2_banks_15_bank_port_2 = (sram_2_ports_cmd_valid && sram_2_ports_cmd_payload_wen[15]);
  assign _zz_sram_3_banks_0_bank_port = sram_3_ports_cmd_payload_wdata[31 : 0];
  assign _zz_sram_3_banks_0_bank_port_1 = sram_3_ports_cmd_payload_wstrb[3 : 0];
  assign _zz_sram_3_banks_0_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[0]);
  assign _zz_sram_3_banks_1_bank_port = sram_3_ports_cmd_payload_wdata[63 : 32];
  assign _zz_sram_3_banks_1_bank_port_1 = sram_3_ports_cmd_payload_wstrb[7 : 4];
  assign _zz_sram_3_banks_1_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[1]);
  assign _zz_sram_3_banks_2_bank_port = sram_3_ports_cmd_payload_wdata[95 : 64];
  assign _zz_sram_3_banks_2_bank_port_1 = sram_3_ports_cmd_payload_wstrb[11 : 8];
  assign _zz_sram_3_banks_2_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[2]);
  assign _zz_sram_3_banks_3_bank_port = sram_3_ports_cmd_payload_wdata[127 : 96];
  assign _zz_sram_3_banks_3_bank_port_1 = sram_3_ports_cmd_payload_wstrb[15 : 12];
  assign _zz_sram_3_banks_3_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[3]);
  assign _zz_sram_3_banks_4_bank_port = sram_3_ports_cmd_payload_wdata[159 : 128];
  assign _zz_sram_3_banks_4_bank_port_1 = sram_3_ports_cmd_payload_wstrb[19 : 16];
  assign _zz_sram_3_banks_4_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[4]);
  assign _zz_sram_3_banks_5_bank_port = sram_3_ports_cmd_payload_wdata[191 : 160];
  assign _zz_sram_3_banks_5_bank_port_1 = sram_3_ports_cmd_payload_wstrb[23 : 20];
  assign _zz_sram_3_banks_5_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[5]);
  assign _zz_sram_3_banks_6_bank_port = sram_3_ports_cmd_payload_wdata[223 : 192];
  assign _zz_sram_3_banks_6_bank_port_1 = sram_3_ports_cmd_payload_wstrb[27 : 24];
  assign _zz_sram_3_banks_6_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[6]);
  assign _zz_sram_3_banks_7_bank_port = sram_3_ports_cmd_payload_wdata[255 : 224];
  assign _zz_sram_3_banks_7_bank_port_1 = sram_3_ports_cmd_payload_wstrb[31 : 28];
  assign _zz_sram_3_banks_7_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[7]);
  assign _zz_sram_3_banks_8_bank_port = sram_3_ports_cmd_payload_wdata[287 : 256];
  assign _zz_sram_3_banks_8_bank_port_1 = sram_3_ports_cmd_payload_wstrb[35 : 32];
  assign _zz_sram_3_banks_8_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[8]);
  assign _zz_sram_3_banks_9_bank_port = sram_3_ports_cmd_payload_wdata[319 : 288];
  assign _zz_sram_3_banks_9_bank_port_1 = sram_3_ports_cmd_payload_wstrb[39 : 36];
  assign _zz_sram_3_banks_9_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[9]);
  assign _zz_sram_3_banks_10_bank_port = sram_3_ports_cmd_payload_wdata[351 : 320];
  assign _zz_sram_3_banks_10_bank_port_1 = sram_3_ports_cmd_payload_wstrb[43 : 40];
  assign _zz_sram_3_banks_10_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[10]);
  assign _zz_sram_3_banks_11_bank_port = sram_3_ports_cmd_payload_wdata[383 : 352];
  assign _zz_sram_3_banks_11_bank_port_1 = sram_3_ports_cmd_payload_wstrb[47 : 44];
  assign _zz_sram_3_banks_11_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[11]);
  assign _zz_sram_3_banks_12_bank_port = sram_3_ports_cmd_payload_wdata[415 : 384];
  assign _zz_sram_3_banks_12_bank_port_1 = sram_3_ports_cmd_payload_wstrb[51 : 48];
  assign _zz_sram_3_banks_12_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[12]);
  assign _zz_sram_3_banks_13_bank_port = sram_3_ports_cmd_payload_wdata[447 : 416];
  assign _zz_sram_3_banks_13_bank_port_1 = sram_3_ports_cmd_payload_wstrb[55 : 52];
  assign _zz_sram_3_banks_13_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[13]);
  assign _zz_sram_3_banks_14_bank_port = sram_3_ports_cmd_payload_wdata[479 : 448];
  assign _zz_sram_3_banks_14_bank_port_1 = sram_3_ports_cmd_payload_wstrb[59 : 56];
  assign _zz_sram_3_banks_14_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[14]);
  assign _zz_sram_3_banks_15_bank_port = sram_3_ports_cmd_payload_wdata[511 : 480];
  assign _zz_sram_3_banks_15_bank_port_1 = sram_3_ports_cmd_payload_wstrb[63 : 60];
  assign _zz_sram_3_banks_15_bank_port_2 = (sram_3_ports_cmd_valid && sram_3_ports_cmd_payload_wen[15]);
  always @(*) begin
    _zz_sram_0_banks_0_bank_port1 = {_zz_sram_0_banks_0_banksymbol_read_3, _zz_sram_0_banks_0_banksymbol_read_2, _zz_sram_0_banks_0_banksymbol_read_1, _zz_sram_0_banks_0_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_0_banks_0_bank_port_1[0] && _zz_sram_0_banks_0_bank_port_2) begin
      sram_0_banks_0_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_0_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_0_bank_port_1[1] && _zz_sram_0_banks_0_bank_port_2) begin
      sram_0_banks_0_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_0_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_0_bank_port_1[2] && _zz_sram_0_banks_0_bank_port_2) begin
      sram_0_banks_0_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_0_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_0_bank_port_1[3] && _zz_sram_0_banks_0_bank_port_2) begin
      sram_0_banks_0_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_0_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_0_banksymbol_read <= sram_0_banks_0_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_0_banksymbol_read_1 <= sram_0_banks_0_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_0_banksymbol_read_2 <= sram_0_banks_0_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_0_banksymbol_read_3 <= sram_0_banks_0_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_0_banks_1_bank_port1 = {_zz_sram_0_banks_1_banksymbol_read_3, _zz_sram_0_banks_1_banksymbol_read_2, _zz_sram_0_banks_1_banksymbol_read_1, _zz_sram_0_banks_1_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_0_banks_1_bank_port_1[0] && _zz_sram_0_banks_1_bank_port_2) begin
      sram_0_banks_1_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_1_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_1_bank_port_1[1] && _zz_sram_0_banks_1_bank_port_2) begin
      sram_0_banks_1_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_1_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_1_bank_port_1[2] && _zz_sram_0_banks_1_bank_port_2) begin
      sram_0_banks_1_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_1_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_1_bank_port_1[3] && _zz_sram_0_banks_1_bank_port_2) begin
      sram_0_banks_1_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_1_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_1_banksymbol_read <= sram_0_banks_1_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_1_banksymbol_read_1 <= sram_0_banks_1_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_1_banksymbol_read_2 <= sram_0_banks_1_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_1_banksymbol_read_3 <= sram_0_banks_1_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_0_banks_2_bank_port1 = {_zz_sram_0_banks_2_banksymbol_read_3, _zz_sram_0_banks_2_banksymbol_read_2, _zz_sram_0_banks_2_banksymbol_read_1, _zz_sram_0_banks_2_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_0_banks_2_bank_port_1[0] && _zz_sram_0_banks_2_bank_port_2) begin
      sram_0_banks_2_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_2_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_2_bank_port_1[1] && _zz_sram_0_banks_2_bank_port_2) begin
      sram_0_banks_2_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_2_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_2_bank_port_1[2] && _zz_sram_0_banks_2_bank_port_2) begin
      sram_0_banks_2_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_2_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_2_bank_port_1[3] && _zz_sram_0_banks_2_bank_port_2) begin
      sram_0_banks_2_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_2_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_2_banksymbol_read <= sram_0_banks_2_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_2_banksymbol_read_1 <= sram_0_banks_2_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_2_banksymbol_read_2 <= sram_0_banks_2_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_2_banksymbol_read_3 <= sram_0_banks_2_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_0_banks_3_bank_port1 = {_zz_sram_0_banks_3_banksymbol_read_3, _zz_sram_0_banks_3_banksymbol_read_2, _zz_sram_0_banks_3_banksymbol_read_1, _zz_sram_0_banks_3_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_0_banks_3_bank_port_1[0] && _zz_sram_0_banks_3_bank_port_2) begin
      sram_0_banks_3_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_3_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_3_bank_port_1[1] && _zz_sram_0_banks_3_bank_port_2) begin
      sram_0_banks_3_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_3_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_3_bank_port_1[2] && _zz_sram_0_banks_3_bank_port_2) begin
      sram_0_banks_3_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_3_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_3_bank_port_1[3] && _zz_sram_0_banks_3_bank_port_2) begin
      sram_0_banks_3_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_3_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_3_banksymbol_read <= sram_0_banks_3_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_3_banksymbol_read_1 <= sram_0_banks_3_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_3_banksymbol_read_2 <= sram_0_banks_3_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_3_banksymbol_read_3 <= sram_0_banks_3_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_0_banks_4_bank_port1 = {_zz_sram_0_banks_4_banksymbol_read_3, _zz_sram_0_banks_4_banksymbol_read_2, _zz_sram_0_banks_4_banksymbol_read_1, _zz_sram_0_banks_4_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_0_banks_4_bank_port_1[0] && _zz_sram_0_banks_4_bank_port_2) begin
      sram_0_banks_4_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_4_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_4_bank_port_1[1] && _zz_sram_0_banks_4_bank_port_2) begin
      sram_0_banks_4_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_4_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_4_bank_port_1[2] && _zz_sram_0_banks_4_bank_port_2) begin
      sram_0_banks_4_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_4_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_4_bank_port_1[3] && _zz_sram_0_banks_4_bank_port_2) begin
      sram_0_banks_4_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_4_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_4_banksymbol_read <= sram_0_banks_4_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_4_banksymbol_read_1 <= sram_0_banks_4_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_4_banksymbol_read_2 <= sram_0_banks_4_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_4_banksymbol_read_3 <= sram_0_banks_4_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_0_banks_5_bank_port1 = {_zz_sram_0_banks_5_banksymbol_read_3, _zz_sram_0_banks_5_banksymbol_read_2, _zz_sram_0_banks_5_banksymbol_read_1, _zz_sram_0_banks_5_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_0_banks_5_bank_port_1[0] && _zz_sram_0_banks_5_bank_port_2) begin
      sram_0_banks_5_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_5_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_5_bank_port_1[1] && _zz_sram_0_banks_5_bank_port_2) begin
      sram_0_banks_5_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_5_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_5_bank_port_1[2] && _zz_sram_0_banks_5_bank_port_2) begin
      sram_0_banks_5_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_5_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_5_bank_port_1[3] && _zz_sram_0_banks_5_bank_port_2) begin
      sram_0_banks_5_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_5_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_5_banksymbol_read <= sram_0_banks_5_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_5_banksymbol_read_1 <= sram_0_banks_5_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_5_banksymbol_read_2 <= sram_0_banks_5_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_5_banksymbol_read_3 <= sram_0_banks_5_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_0_banks_6_bank_port1 = {_zz_sram_0_banks_6_banksymbol_read_3, _zz_sram_0_banks_6_banksymbol_read_2, _zz_sram_0_banks_6_banksymbol_read_1, _zz_sram_0_banks_6_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_0_banks_6_bank_port_1[0] && _zz_sram_0_banks_6_bank_port_2) begin
      sram_0_banks_6_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_6_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_6_bank_port_1[1] && _zz_sram_0_banks_6_bank_port_2) begin
      sram_0_banks_6_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_6_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_6_bank_port_1[2] && _zz_sram_0_banks_6_bank_port_2) begin
      sram_0_banks_6_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_6_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_6_bank_port_1[3] && _zz_sram_0_banks_6_bank_port_2) begin
      sram_0_banks_6_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_6_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_6_banksymbol_read <= sram_0_banks_6_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_6_banksymbol_read_1 <= sram_0_banks_6_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_6_banksymbol_read_2 <= sram_0_banks_6_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_6_banksymbol_read_3 <= sram_0_banks_6_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_0_banks_7_bank_port1 = {_zz_sram_0_banks_7_banksymbol_read_3, _zz_sram_0_banks_7_banksymbol_read_2, _zz_sram_0_banks_7_banksymbol_read_1, _zz_sram_0_banks_7_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_0_banks_7_bank_port_1[0] && _zz_sram_0_banks_7_bank_port_2) begin
      sram_0_banks_7_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_7_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_7_bank_port_1[1] && _zz_sram_0_banks_7_bank_port_2) begin
      sram_0_banks_7_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_7_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_7_bank_port_1[2] && _zz_sram_0_banks_7_bank_port_2) begin
      sram_0_banks_7_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_7_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_7_bank_port_1[3] && _zz_sram_0_banks_7_bank_port_2) begin
      sram_0_banks_7_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_7_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_7_banksymbol_read <= sram_0_banks_7_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_7_banksymbol_read_1 <= sram_0_banks_7_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_7_banksymbol_read_2 <= sram_0_banks_7_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_7_banksymbol_read_3 <= sram_0_banks_7_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_0_banks_8_bank_port1 = {_zz_sram_0_banks_8_banksymbol_read_3, _zz_sram_0_banks_8_banksymbol_read_2, _zz_sram_0_banks_8_banksymbol_read_1, _zz_sram_0_banks_8_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_0_banks_8_bank_port_1[0] && _zz_sram_0_banks_8_bank_port_2) begin
      sram_0_banks_8_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_8_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_8_bank_port_1[1] && _zz_sram_0_banks_8_bank_port_2) begin
      sram_0_banks_8_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_8_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_8_bank_port_1[2] && _zz_sram_0_banks_8_bank_port_2) begin
      sram_0_banks_8_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_8_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_8_bank_port_1[3] && _zz_sram_0_banks_8_bank_port_2) begin
      sram_0_banks_8_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_8_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_8_banksymbol_read <= sram_0_banks_8_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_8_banksymbol_read_1 <= sram_0_banks_8_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_8_banksymbol_read_2 <= sram_0_banks_8_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_8_banksymbol_read_3 <= sram_0_banks_8_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_0_banks_9_bank_port1 = {_zz_sram_0_banks_9_banksymbol_read_3, _zz_sram_0_banks_9_banksymbol_read_2, _zz_sram_0_banks_9_banksymbol_read_1, _zz_sram_0_banks_9_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_0_banks_9_bank_port_1[0] && _zz_sram_0_banks_9_bank_port_2) begin
      sram_0_banks_9_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_9_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_9_bank_port_1[1] && _zz_sram_0_banks_9_bank_port_2) begin
      sram_0_banks_9_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_9_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_9_bank_port_1[2] && _zz_sram_0_banks_9_bank_port_2) begin
      sram_0_banks_9_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_9_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_9_bank_port_1[3] && _zz_sram_0_banks_9_bank_port_2) begin
      sram_0_banks_9_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_9_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_9_banksymbol_read <= sram_0_banks_9_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_9_banksymbol_read_1 <= sram_0_banks_9_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_9_banksymbol_read_2 <= sram_0_banks_9_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_9_banksymbol_read_3 <= sram_0_banks_9_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_0_banks_10_bank_port1 = {_zz_sram_0_banks_10_banksymbol_read_3, _zz_sram_0_banks_10_banksymbol_read_2, _zz_sram_0_banks_10_banksymbol_read_1, _zz_sram_0_banks_10_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_0_banks_10_bank_port_1[0] && _zz_sram_0_banks_10_bank_port_2) begin
      sram_0_banks_10_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_10_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_10_bank_port_1[1] && _zz_sram_0_banks_10_bank_port_2) begin
      sram_0_banks_10_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_10_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_10_bank_port_1[2] && _zz_sram_0_banks_10_bank_port_2) begin
      sram_0_banks_10_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_10_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_10_bank_port_1[3] && _zz_sram_0_banks_10_bank_port_2) begin
      sram_0_banks_10_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_10_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_10_banksymbol_read <= sram_0_banks_10_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_10_banksymbol_read_1 <= sram_0_banks_10_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_10_banksymbol_read_2 <= sram_0_banks_10_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_10_banksymbol_read_3 <= sram_0_banks_10_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_0_banks_11_bank_port1 = {_zz_sram_0_banks_11_banksymbol_read_3, _zz_sram_0_banks_11_banksymbol_read_2, _zz_sram_0_banks_11_banksymbol_read_1, _zz_sram_0_banks_11_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_0_banks_11_bank_port_1[0] && _zz_sram_0_banks_11_bank_port_2) begin
      sram_0_banks_11_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_11_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_11_bank_port_1[1] && _zz_sram_0_banks_11_bank_port_2) begin
      sram_0_banks_11_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_11_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_11_bank_port_1[2] && _zz_sram_0_banks_11_bank_port_2) begin
      sram_0_banks_11_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_11_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_11_bank_port_1[3] && _zz_sram_0_banks_11_bank_port_2) begin
      sram_0_banks_11_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_11_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_11_banksymbol_read <= sram_0_banks_11_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_11_banksymbol_read_1 <= sram_0_banks_11_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_11_banksymbol_read_2 <= sram_0_banks_11_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_11_banksymbol_read_3 <= sram_0_banks_11_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_0_banks_12_bank_port1 = {_zz_sram_0_banks_12_banksymbol_read_3, _zz_sram_0_banks_12_banksymbol_read_2, _zz_sram_0_banks_12_banksymbol_read_1, _zz_sram_0_banks_12_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_0_banks_12_bank_port_1[0] && _zz_sram_0_banks_12_bank_port_2) begin
      sram_0_banks_12_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_12_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_12_bank_port_1[1] && _zz_sram_0_banks_12_bank_port_2) begin
      sram_0_banks_12_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_12_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_12_bank_port_1[2] && _zz_sram_0_banks_12_bank_port_2) begin
      sram_0_banks_12_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_12_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_12_bank_port_1[3] && _zz_sram_0_banks_12_bank_port_2) begin
      sram_0_banks_12_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_12_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_12_banksymbol_read <= sram_0_banks_12_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_12_banksymbol_read_1 <= sram_0_banks_12_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_12_banksymbol_read_2 <= sram_0_banks_12_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_12_banksymbol_read_3 <= sram_0_banks_12_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_0_banks_13_bank_port1 = {_zz_sram_0_banks_13_banksymbol_read_3, _zz_sram_0_banks_13_banksymbol_read_2, _zz_sram_0_banks_13_banksymbol_read_1, _zz_sram_0_banks_13_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_0_banks_13_bank_port_1[0] && _zz_sram_0_banks_13_bank_port_2) begin
      sram_0_banks_13_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_13_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_13_bank_port_1[1] && _zz_sram_0_banks_13_bank_port_2) begin
      sram_0_banks_13_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_13_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_13_bank_port_1[2] && _zz_sram_0_banks_13_bank_port_2) begin
      sram_0_banks_13_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_13_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_13_bank_port_1[3] && _zz_sram_0_banks_13_bank_port_2) begin
      sram_0_banks_13_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_13_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_13_banksymbol_read <= sram_0_banks_13_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_13_banksymbol_read_1 <= sram_0_banks_13_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_13_banksymbol_read_2 <= sram_0_banks_13_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_13_banksymbol_read_3 <= sram_0_banks_13_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_0_banks_14_bank_port1 = {_zz_sram_0_banks_14_banksymbol_read_3, _zz_sram_0_banks_14_banksymbol_read_2, _zz_sram_0_banks_14_banksymbol_read_1, _zz_sram_0_banks_14_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_0_banks_14_bank_port_1[0] && _zz_sram_0_banks_14_bank_port_2) begin
      sram_0_banks_14_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_14_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_14_bank_port_1[1] && _zz_sram_0_banks_14_bank_port_2) begin
      sram_0_banks_14_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_14_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_14_bank_port_1[2] && _zz_sram_0_banks_14_bank_port_2) begin
      sram_0_banks_14_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_14_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_14_bank_port_1[3] && _zz_sram_0_banks_14_bank_port_2) begin
      sram_0_banks_14_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_14_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_14_banksymbol_read <= sram_0_banks_14_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_14_banksymbol_read_1 <= sram_0_banks_14_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_14_banksymbol_read_2 <= sram_0_banks_14_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_14_banksymbol_read_3 <= sram_0_banks_14_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_0_banks_15_bank_port1 = {_zz_sram_0_banks_15_banksymbol_read_3, _zz_sram_0_banks_15_banksymbol_read_2, _zz_sram_0_banks_15_banksymbol_read_1, _zz_sram_0_banks_15_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_0_banks_15_bank_port_1[0] && _zz_sram_0_banks_15_bank_port_2) begin
      sram_0_banks_15_bank_symbol0[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_15_bank_port[7 : 0];
    end
    if(_zz_sram_0_banks_15_bank_port_1[1] && _zz_sram_0_banks_15_bank_port_2) begin
      sram_0_banks_15_bank_symbol1[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_15_bank_port[15 : 8];
    end
    if(_zz_sram_0_banks_15_bank_port_1[2] && _zz_sram_0_banks_15_bank_port_2) begin
      sram_0_banks_15_bank_symbol2[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_15_bank_port[23 : 16];
    end
    if(_zz_sram_0_banks_15_bank_port_1[3] && _zz_sram_0_banks_15_bank_port_2) begin
      sram_0_banks_15_bank_symbol3[sram_0_ports_cmd_payload_addr] <= _zz_sram_0_banks_15_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_0_ports_cmd_valid) begin
      _zz_sram_0_banks_15_banksymbol_read <= sram_0_banks_15_bank_symbol0[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_15_banksymbol_read_1 <= sram_0_banks_15_bank_symbol1[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_15_banksymbol_read_2 <= sram_0_banks_15_bank_symbol2[sram_0_ports_cmd_payload_addr];
      _zz_sram_0_banks_15_banksymbol_read_3 <= sram_0_banks_15_bank_symbol3[sram_0_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_0_bank_port1 = {_zz_sram_1_banks_0_banksymbol_read_3, _zz_sram_1_banks_0_banksymbol_read_2, _zz_sram_1_banks_0_banksymbol_read_1, _zz_sram_1_banks_0_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_1_banks_0_bank_port_1[0] && _zz_sram_1_banks_0_bank_port_2) begin
      sram_1_banks_0_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_0_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_0_bank_port_1[1] && _zz_sram_1_banks_0_bank_port_2) begin
      sram_1_banks_0_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_0_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_0_bank_port_1[2] && _zz_sram_1_banks_0_bank_port_2) begin
      sram_1_banks_0_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_0_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_0_bank_port_1[3] && _zz_sram_1_banks_0_bank_port_2) begin
      sram_1_banks_0_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_0_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_0_banksymbol_read <= sram_1_banks_0_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_0_banksymbol_read_1 <= sram_1_banks_0_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_0_banksymbol_read_2 <= sram_1_banks_0_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_0_banksymbol_read_3 <= sram_1_banks_0_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_1_bank_port1 = {_zz_sram_1_banks_1_banksymbol_read_3, _zz_sram_1_banks_1_banksymbol_read_2, _zz_sram_1_banks_1_banksymbol_read_1, _zz_sram_1_banks_1_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_1_banks_1_bank_port_1[0] && _zz_sram_1_banks_1_bank_port_2) begin
      sram_1_banks_1_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_1_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_1_bank_port_1[1] && _zz_sram_1_banks_1_bank_port_2) begin
      sram_1_banks_1_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_1_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_1_bank_port_1[2] && _zz_sram_1_banks_1_bank_port_2) begin
      sram_1_banks_1_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_1_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_1_bank_port_1[3] && _zz_sram_1_banks_1_bank_port_2) begin
      sram_1_banks_1_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_1_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_1_banksymbol_read <= sram_1_banks_1_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_1_banksymbol_read_1 <= sram_1_banks_1_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_1_banksymbol_read_2 <= sram_1_banks_1_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_1_banksymbol_read_3 <= sram_1_banks_1_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_2_bank_port1 = {_zz_sram_1_banks_2_banksymbol_read_3, _zz_sram_1_banks_2_banksymbol_read_2, _zz_sram_1_banks_2_banksymbol_read_1, _zz_sram_1_banks_2_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_1_banks_2_bank_port_1[0] && _zz_sram_1_banks_2_bank_port_2) begin
      sram_1_banks_2_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_2_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_2_bank_port_1[1] && _zz_sram_1_banks_2_bank_port_2) begin
      sram_1_banks_2_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_2_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_2_bank_port_1[2] && _zz_sram_1_banks_2_bank_port_2) begin
      sram_1_banks_2_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_2_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_2_bank_port_1[3] && _zz_sram_1_banks_2_bank_port_2) begin
      sram_1_banks_2_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_2_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_2_banksymbol_read <= sram_1_banks_2_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_2_banksymbol_read_1 <= sram_1_banks_2_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_2_banksymbol_read_2 <= sram_1_banks_2_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_2_banksymbol_read_3 <= sram_1_banks_2_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_3_bank_port1 = {_zz_sram_1_banks_3_banksymbol_read_3, _zz_sram_1_banks_3_banksymbol_read_2, _zz_sram_1_banks_3_banksymbol_read_1, _zz_sram_1_banks_3_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_1_banks_3_bank_port_1[0] && _zz_sram_1_banks_3_bank_port_2) begin
      sram_1_banks_3_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_3_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_3_bank_port_1[1] && _zz_sram_1_banks_3_bank_port_2) begin
      sram_1_banks_3_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_3_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_3_bank_port_1[2] && _zz_sram_1_banks_3_bank_port_2) begin
      sram_1_banks_3_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_3_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_3_bank_port_1[3] && _zz_sram_1_banks_3_bank_port_2) begin
      sram_1_banks_3_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_3_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_3_banksymbol_read <= sram_1_banks_3_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_3_banksymbol_read_1 <= sram_1_banks_3_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_3_banksymbol_read_2 <= sram_1_banks_3_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_3_banksymbol_read_3 <= sram_1_banks_3_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_4_bank_port1 = {_zz_sram_1_banks_4_banksymbol_read_3, _zz_sram_1_banks_4_banksymbol_read_2, _zz_sram_1_banks_4_banksymbol_read_1, _zz_sram_1_banks_4_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_1_banks_4_bank_port_1[0] && _zz_sram_1_banks_4_bank_port_2) begin
      sram_1_banks_4_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_4_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_4_bank_port_1[1] && _zz_sram_1_banks_4_bank_port_2) begin
      sram_1_banks_4_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_4_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_4_bank_port_1[2] && _zz_sram_1_banks_4_bank_port_2) begin
      sram_1_banks_4_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_4_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_4_bank_port_1[3] && _zz_sram_1_banks_4_bank_port_2) begin
      sram_1_banks_4_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_4_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_4_banksymbol_read <= sram_1_banks_4_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_4_banksymbol_read_1 <= sram_1_banks_4_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_4_banksymbol_read_2 <= sram_1_banks_4_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_4_banksymbol_read_3 <= sram_1_banks_4_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_5_bank_port1 = {_zz_sram_1_banks_5_banksymbol_read_3, _zz_sram_1_banks_5_banksymbol_read_2, _zz_sram_1_banks_5_banksymbol_read_1, _zz_sram_1_banks_5_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_1_banks_5_bank_port_1[0] && _zz_sram_1_banks_5_bank_port_2) begin
      sram_1_banks_5_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_5_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_5_bank_port_1[1] && _zz_sram_1_banks_5_bank_port_2) begin
      sram_1_banks_5_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_5_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_5_bank_port_1[2] && _zz_sram_1_banks_5_bank_port_2) begin
      sram_1_banks_5_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_5_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_5_bank_port_1[3] && _zz_sram_1_banks_5_bank_port_2) begin
      sram_1_banks_5_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_5_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_5_banksymbol_read <= sram_1_banks_5_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_5_banksymbol_read_1 <= sram_1_banks_5_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_5_banksymbol_read_2 <= sram_1_banks_5_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_5_banksymbol_read_3 <= sram_1_banks_5_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_6_bank_port1 = {_zz_sram_1_banks_6_banksymbol_read_3, _zz_sram_1_banks_6_banksymbol_read_2, _zz_sram_1_banks_6_banksymbol_read_1, _zz_sram_1_banks_6_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_1_banks_6_bank_port_1[0] && _zz_sram_1_banks_6_bank_port_2) begin
      sram_1_banks_6_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_6_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_6_bank_port_1[1] && _zz_sram_1_banks_6_bank_port_2) begin
      sram_1_banks_6_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_6_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_6_bank_port_1[2] && _zz_sram_1_banks_6_bank_port_2) begin
      sram_1_banks_6_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_6_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_6_bank_port_1[3] && _zz_sram_1_banks_6_bank_port_2) begin
      sram_1_banks_6_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_6_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_6_banksymbol_read <= sram_1_banks_6_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_6_banksymbol_read_1 <= sram_1_banks_6_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_6_banksymbol_read_2 <= sram_1_banks_6_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_6_banksymbol_read_3 <= sram_1_banks_6_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_7_bank_port1 = {_zz_sram_1_banks_7_banksymbol_read_3, _zz_sram_1_banks_7_banksymbol_read_2, _zz_sram_1_banks_7_banksymbol_read_1, _zz_sram_1_banks_7_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_1_banks_7_bank_port_1[0] && _zz_sram_1_banks_7_bank_port_2) begin
      sram_1_banks_7_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_7_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_7_bank_port_1[1] && _zz_sram_1_banks_7_bank_port_2) begin
      sram_1_banks_7_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_7_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_7_bank_port_1[2] && _zz_sram_1_banks_7_bank_port_2) begin
      sram_1_banks_7_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_7_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_7_bank_port_1[3] && _zz_sram_1_banks_7_bank_port_2) begin
      sram_1_banks_7_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_7_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_7_banksymbol_read <= sram_1_banks_7_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_7_banksymbol_read_1 <= sram_1_banks_7_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_7_banksymbol_read_2 <= sram_1_banks_7_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_7_banksymbol_read_3 <= sram_1_banks_7_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_8_bank_port1 = {_zz_sram_1_banks_8_banksymbol_read_3, _zz_sram_1_banks_8_banksymbol_read_2, _zz_sram_1_banks_8_banksymbol_read_1, _zz_sram_1_banks_8_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_1_banks_8_bank_port_1[0] && _zz_sram_1_banks_8_bank_port_2) begin
      sram_1_banks_8_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_8_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_8_bank_port_1[1] && _zz_sram_1_banks_8_bank_port_2) begin
      sram_1_banks_8_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_8_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_8_bank_port_1[2] && _zz_sram_1_banks_8_bank_port_2) begin
      sram_1_banks_8_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_8_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_8_bank_port_1[3] && _zz_sram_1_banks_8_bank_port_2) begin
      sram_1_banks_8_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_8_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_8_banksymbol_read <= sram_1_banks_8_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_8_banksymbol_read_1 <= sram_1_banks_8_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_8_banksymbol_read_2 <= sram_1_banks_8_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_8_banksymbol_read_3 <= sram_1_banks_8_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_9_bank_port1 = {_zz_sram_1_banks_9_banksymbol_read_3, _zz_sram_1_banks_9_banksymbol_read_2, _zz_sram_1_banks_9_banksymbol_read_1, _zz_sram_1_banks_9_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_1_banks_9_bank_port_1[0] && _zz_sram_1_banks_9_bank_port_2) begin
      sram_1_banks_9_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_9_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_9_bank_port_1[1] && _zz_sram_1_banks_9_bank_port_2) begin
      sram_1_banks_9_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_9_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_9_bank_port_1[2] && _zz_sram_1_banks_9_bank_port_2) begin
      sram_1_banks_9_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_9_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_9_bank_port_1[3] && _zz_sram_1_banks_9_bank_port_2) begin
      sram_1_banks_9_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_9_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_9_banksymbol_read <= sram_1_banks_9_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_9_banksymbol_read_1 <= sram_1_banks_9_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_9_banksymbol_read_2 <= sram_1_banks_9_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_9_banksymbol_read_3 <= sram_1_banks_9_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_10_bank_port1 = {_zz_sram_1_banks_10_banksymbol_read_3, _zz_sram_1_banks_10_banksymbol_read_2, _zz_sram_1_banks_10_banksymbol_read_1, _zz_sram_1_banks_10_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_1_banks_10_bank_port_1[0] && _zz_sram_1_banks_10_bank_port_2) begin
      sram_1_banks_10_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_10_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_10_bank_port_1[1] && _zz_sram_1_banks_10_bank_port_2) begin
      sram_1_banks_10_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_10_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_10_bank_port_1[2] && _zz_sram_1_banks_10_bank_port_2) begin
      sram_1_banks_10_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_10_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_10_bank_port_1[3] && _zz_sram_1_banks_10_bank_port_2) begin
      sram_1_banks_10_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_10_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_10_banksymbol_read <= sram_1_banks_10_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_10_banksymbol_read_1 <= sram_1_banks_10_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_10_banksymbol_read_2 <= sram_1_banks_10_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_10_banksymbol_read_3 <= sram_1_banks_10_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_11_bank_port1 = {_zz_sram_1_banks_11_banksymbol_read_3, _zz_sram_1_banks_11_banksymbol_read_2, _zz_sram_1_banks_11_banksymbol_read_1, _zz_sram_1_banks_11_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_1_banks_11_bank_port_1[0] && _zz_sram_1_banks_11_bank_port_2) begin
      sram_1_banks_11_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_11_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_11_bank_port_1[1] && _zz_sram_1_banks_11_bank_port_2) begin
      sram_1_banks_11_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_11_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_11_bank_port_1[2] && _zz_sram_1_banks_11_bank_port_2) begin
      sram_1_banks_11_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_11_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_11_bank_port_1[3] && _zz_sram_1_banks_11_bank_port_2) begin
      sram_1_banks_11_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_11_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_11_banksymbol_read <= sram_1_banks_11_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_11_banksymbol_read_1 <= sram_1_banks_11_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_11_banksymbol_read_2 <= sram_1_banks_11_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_11_banksymbol_read_3 <= sram_1_banks_11_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_12_bank_port1 = {_zz_sram_1_banks_12_banksymbol_read_3, _zz_sram_1_banks_12_banksymbol_read_2, _zz_sram_1_banks_12_banksymbol_read_1, _zz_sram_1_banks_12_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_1_banks_12_bank_port_1[0] && _zz_sram_1_banks_12_bank_port_2) begin
      sram_1_banks_12_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_12_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_12_bank_port_1[1] && _zz_sram_1_banks_12_bank_port_2) begin
      sram_1_banks_12_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_12_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_12_bank_port_1[2] && _zz_sram_1_banks_12_bank_port_2) begin
      sram_1_banks_12_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_12_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_12_bank_port_1[3] && _zz_sram_1_banks_12_bank_port_2) begin
      sram_1_banks_12_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_12_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_12_banksymbol_read <= sram_1_banks_12_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_12_banksymbol_read_1 <= sram_1_banks_12_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_12_banksymbol_read_2 <= sram_1_banks_12_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_12_banksymbol_read_3 <= sram_1_banks_12_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_13_bank_port1 = {_zz_sram_1_banks_13_banksymbol_read_3, _zz_sram_1_banks_13_banksymbol_read_2, _zz_sram_1_banks_13_banksymbol_read_1, _zz_sram_1_banks_13_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_1_banks_13_bank_port_1[0] && _zz_sram_1_banks_13_bank_port_2) begin
      sram_1_banks_13_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_13_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_13_bank_port_1[1] && _zz_sram_1_banks_13_bank_port_2) begin
      sram_1_banks_13_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_13_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_13_bank_port_1[2] && _zz_sram_1_banks_13_bank_port_2) begin
      sram_1_banks_13_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_13_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_13_bank_port_1[3] && _zz_sram_1_banks_13_bank_port_2) begin
      sram_1_banks_13_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_13_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_13_banksymbol_read <= sram_1_banks_13_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_13_banksymbol_read_1 <= sram_1_banks_13_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_13_banksymbol_read_2 <= sram_1_banks_13_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_13_banksymbol_read_3 <= sram_1_banks_13_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_14_bank_port1 = {_zz_sram_1_banks_14_banksymbol_read_3, _zz_sram_1_banks_14_banksymbol_read_2, _zz_sram_1_banks_14_banksymbol_read_1, _zz_sram_1_banks_14_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_1_banks_14_bank_port_1[0] && _zz_sram_1_banks_14_bank_port_2) begin
      sram_1_banks_14_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_14_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_14_bank_port_1[1] && _zz_sram_1_banks_14_bank_port_2) begin
      sram_1_banks_14_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_14_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_14_bank_port_1[2] && _zz_sram_1_banks_14_bank_port_2) begin
      sram_1_banks_14_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_14_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_14_bank_port_1[3] && _zz_sram_1_banks_14_bank_port_2) begin
      sram_1_banks_14_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_14_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_14_banksymbol_read <= sram_1_banks_14_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_14_banksymbol_read_1 <= sram_1_banks_14_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_14_banksymbol_read_2 <= sram_1_banks_14_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_14_banksymbol_read_3 <= sram_1_banks_14_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_1_banks_15_bank_port1 = {_zz_sram_1_banks_15_banksymbol_read_3, _zz_sram_1_banks_15_banksymbol_read_2, _zz_sram_1_banks_15_banksymbol_read_1, _zz_sram_1_banks_15_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_1_banks_15_bank_port_1[0] && _zz_sram_1_banks_15_bank_port_2) begin
      sram_1_banks_15_bank_symbol0[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_15_bank_port[7 : 0];
    end
    if(_zz_sram_1_banks_15_bank_port_1[1] && _zz_sram_1_banks_15_bank_port_2) begin
      sram_1_banks_15_bank_symbol1[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_15_bank_port[15 : 8];
    end
    if(_zz_sram_1_banks_15_bank_port_1[2] && _zz_sram_1_banks_15_bank_port_2) begin
      sram_1_banks_15_bank_symbol2[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_15_bank_port[23 : 16];
    end
    if(_zz_sram_1_banks_15_bank_port_1[3] && _zz_sram_1_banks_15_bank_port_2) begin
      sram_1_banks_15_bank_symbol3[sram_1_ports_cmd_payload_addr] <= _zz_sram_1_banks_15_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_1_ports_cmd_valid) begin
      _zz_sram_1_banks_15_banksymbol_read <= sram_1_banks_15_bank_symbol0[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_15_banksymbol_read_1 <= sram_1_banks_15_bank_symbol1[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_15_banksymbol_read_2 <= sram_1_banks_15_bank_symbol2[sram_1_ports_cmd_payload_addr];
      _zz_sram_1_banks_15_banksymbol_read_3 <= sram_1_banks_15_bank_symbol3[sram_1_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_0_bank_port1 = {_zz_sram_2_banks_0_banksymbol_read_3, _zz_sram_2_banks_0_banksymbol_read_2, _zz_sram_2_banks_0_banksymbol_read_1, _zz_sram_2_banks_0_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_2_banks_0_bank_port_1[0] && _zz_sram_2_banks_0_bank_port_2) begin
      sram_2_banks_0_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_0_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_0_bank_port_1[1] && _zz_sram_2_banks_0_bank_port_2) begin
      sram_2_banks_0_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_0_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_0_bank_port_1[2] && _zz_sram_2_banks_0_bank_port_2) begin
      sram_2_banks_0_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_0_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_0_bank_port_1[3] && _zz_sram_2_banks_0_bank_port_2) begin
      sram_2_banks_0_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_0_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_0_banksymbol_read <= sram_2_banks_0_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_0_banksymbol_read_1 <= sram_2_banks_0_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_0_banksymbol_read_2 <= sram_2_banks_0_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_0_banksymbol_read_3 <= sram_2_banks_0_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_1_bank_port1 = {_zz_sram_2_banks_1_banksymbol_read_3, _zz_sram_2_banks_1_banksymbol_read_2, _zz_sram_2_banks_1_banksymbol_read_1, _zz_sram_2_banks_1_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_2_banks_1_bank_port_1[0] && _zz_sram_2_banks_1_bank_port_2) begin
      sram_2_banks_1_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_1_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_1_bank_port_1[1] && _zz_sram_2_banks_1_bank_port_2) begin
      sram_2_banks_1_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_1_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_1_bank_port_1[2] && _zz_sram_2_banks_1_bank_port_2) begin
      sram_2_banks_1_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_1_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_1_bank_port_1[3] && _zz_sram_2_banks_1_bank_port_2) begin
      sram_2_banks_1_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_1_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_1_banksymbol_read <= sram_2_banks_1_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_1_banksymbol_read_1 <= sram_2_banks_1_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_1_banksymbol_read_2 <= sram_2_banks_1_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_1_banksymbol_read_3 <= sram_2_banks_1_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_2_bank_port1 = {_zz_sram_2_banks_2_banksymbol_read_3, _zz_sram_2_banks_2_banksymbol_read_2, _zz_sram_2_banks_2_banksymbol_read_1, _zz_sram_2_banks_2_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_2_banks_2_bank_port_1[0] && _zz_sram_2_banks_2_bank_port_2) begin
      sram_2_banks_2_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_2_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_2_bank_port_1[1] && _zz_sram_2_banks_2_bank_port_2) begin
      sram_2_banks_2_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_2_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_2_bank_port_1[2] && _zz_sram_2_banks_2_bank_port_2) begin
      sram_2_banks_2_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_2_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_2_bank_port_1[3] && _zz_sram_2_banks_2_bank_port_2) begin
      sram_2_banks_2_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_2_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_2_banksymbol_read <= sram_2_banks_2_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_2_banksymbol_read_1 <= sram_2_banks_2_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_2_banksymbol_read_2 <= sram_2_banks_2_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_2_banksymbol_read_3 <= sram_2_banks_2_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_3_bank_port1 = {_zz_sram_2_banks_3_banksymbol_read_3, _zz_sram_2_banks_3_banksymbol_read_2, _zz_sram_2_banks_3_banksymbol_read_1, _zz_sram_2_banks_3_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_2_banks_3_bank_port_1[0] && _zz_sram_2_banks_3_bank_port_2) begin
      sram_2_banks_3_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_3_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_3_bank_port_1[1] && _zz_sram_2_banks_3_bank_port_2) begin
      sram_2_banks_3_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_3_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_3_bank_port_1[2] && _zz_sram_2_banks_3_bank_port_2) begin
      sram_2_banks_3_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_3_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_3_bank_port_1[3] && _zz_sram_2_banks_3_bank_port_2) begin
      sram_2_banks_3_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_3_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_3_banksymbol_read <= sram_2_banks_3_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_3_banksymbol_read_1 <= sram_2_banks_3_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_3_banksymbol_read_2 <= sram_2_banks_3_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_3_banksymbol_read_3 <= sram_2_banks_3_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_4_bank_port1 = {_zz_sram_2_banks_4_banksymbol_read_3, _zz_sram_2_banks_4_banksymbol_read_2, _zz_sram_2_banks_4_banksymbol_read_1, _zz_sram_2_banks_4_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_2_banks_4_bank_port_1[0] && _zz_sram_2_banks_4_bank_port_2) begin
      sram_2_banks_4_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_4_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_4_bank_port_1[1] && _zz_sram_2_banks_4_bank_port_2) begin
      sram_2_banks_4_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_4_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_4_bank_port_1[2] && _zz_sram_2_banks_4_bank_port_2) begin
      sram_2_banks_4_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_4_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_4_bank_port_1[3] && _zz_sram_2_banks_4_bank_port_2) begin
      sram_2_banks_4_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_4_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_4_banksymbol_read <= sram_2_banks_4_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_4_banksymbol_read_1 <= sram_2_banks_4_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_4_banksymbol_read_2 <= sram_2_banks_4_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_4_banksymbol_read_3 <= sram_2_banks_4_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_5_bank_port1 = {_zz_sram_2_banks_5_banksymbol_read_3, _zz_sram_2_banks_5_banksymbol_read_2, _zz_sram_2_banks_5_banksymbol_read_1, _zz_sram_2_banks_5_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_2_banks_5_bank_port_1[0] && _zz_sram_2_banks_5_bank_port_2) begin
      sram_2_banks_5_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_5_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_5_bank_port_1[1] && _zz_sram_2_banks_5_bank_port_2) begin
      sram_2_banks_5_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_5_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_5_bank_port_1[2] && _zz_sram_2_banks_5_bank_port_2) begin
      sram_2_banks_5_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_5_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_5_bank_port_1[3] && _zz_sram_2_banks_5_bank_port_2) begin
      sram_2_banks_5_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_5_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_5_banksymbol_read <= sram_2_banks_5_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_5_banksymbol_read_1 <= sram_2_banks_5_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_5_banksymbol_read_2 <= sram_2_banks_5_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_5_banksymbol_read_3 <= sram_2_banks_5_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_6_bank_port1 = {_zz_sram_2_banks_6_banksymbol_read_3, _zz_sram_2_banks_6_banksymbol_read_2, _zz_sram_2_banks_6_banksymbol_read_1, _zz_sram_2_banks_6_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_2_banks_6_bank_port_1[0] && _zz_sram_2_banks_6_bank_port_2) begin
      sram_2_banks_6_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_6_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_6_bank_port_1[1] && _zz_sram_2_banks_6_bank_port_2) begin
      sram_2_banks_6_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_6_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_6_bank_port_1[2] && _zz_sram_2_banks_6_bank_port_2) begin
      sram_2_banks_6_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_6_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_6_bank_port_1[3] && _zz_sram_2_banks_6_bank_port_2) begin
      sram_2_banks_6_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_6_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_6_banksymbol_read <= sram_2_banks_6_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_6_banksymbol_read_1 <= sram_2_banks_6_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_6_banksymbol_read_2 <= sram_2_banks_6_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_6_banksymbol_read_3 <= sram_2_banks_6_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_7_bank_port1 = {_zz_sram_2_banks_7_banksymbol_read_3, _zz_sram_2_banks_7_banksymbol_read_2, _zz_sram_2_banks_7_banksymbol_read_1, _zz_sram_2_banks_7_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_2_banks_7_bank_port_1[0] && _zz_sram_2_banks_7_bank_port_2) begin
      sram_2_banks_7_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_7_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_7_bank_port_1[1] && _zz_sram_2_banks_7_bank_port_2) begin
      sram_2_banks_7_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_7_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_7_bank_port_1[2] && _zz_sram_2_banks_7_bank_port_2) begin
      sram_2_banks_7_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_7_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_7_bank_port_1[3] && _zz_sram_2_banks_7_bank_port_2) begin
      sram_2_banks_7_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_7_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_7_banksymbol_read <= sram_2_banks_7_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_7_banksymbol_read_1 <= sram_2_banks_7_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_7_banksymbol_read_2 <= sram_2_banks_7_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_7_banksymbol_read_3 <= sram_2_banks_7_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_8_bank_port1 = {_zz_sram_2_banks_8_banksymbol_read_3, _zz_sram_2_banks_8_banksymbol_read_2, _zz_sram_2_banks_8_banksymbol_read_1, _zz_sram_2_banks_8_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_2_banks_8_bank_port_1[0] && _zz_sram_2_banks_8_bank_port_2) begin
      sram_2_banks_8_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_8_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_8_bank_port_1[1] && _zz_sram_2_banks_8_bank_port_2) begin
      sram_2_banks_8_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_8_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_8_bank_port_1[2] && _zz_sram_2_banks_8_bank_port_2) begin
      sram_2_banks_8_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_8_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_8_bank_port_1[3] && _zz_sram_2_banks_8_bank_port_2) begin
      sram_2_banks_8_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_8_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_8_banksymbol_read <= sram_2_banks_8_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_8_banksymbol_read_1 <= sram_2_banks_8_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_8_banksymbol_read_2 <= sram_2_banks_8_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_8_banksymbol_read_3 <= sram_2_banks_8_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_9_bank_port1 = {_zz_sram_2_banks_9_banksymbol_read_3, _zz_sram_2_banks_9_banksymbol_read_2, _zz_sram_2_banks_9_banksymbol_read_1, _zz_sram_2_banks_9_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_2_banks_9_bank_port_1[0] && _zz_sram_2_banks_9_bank_port_2) begin
      sram_2_banks_9_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_9_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_9_bank_port_1[1] && _zz_sram_2_banks_9_bank_port_2) begin
      sram_2_banks_9_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_9_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_9_bank_port_1[2] && _zz_sram_2_banks_9_bank_port_2) begin
      sram_2_banks_9_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_9_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_9_bank_port_1[3] && _zz_sram_2_banks_9_bank_port_2) begin
      sram_2_banks_9_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_9_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_9_banksymbol_read <= sram_2_banks_9_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_9_banksymbol_read_1 <= sram_2_banks_9_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_9_banksymbol_read_2 <= sram_2_banks_9_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_9_banksymbol_read_3 <= sram_2_banks_9_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_10_bank_port1 = {_zz_sram_2_banks_10_banksymbol_read_3, _zz_sram_2_banks_10_banksymbol_read_2, _zz_sram_2_banks_10_banksymbol_read_1, _zz_sram_2_banks_10_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_2_banks_10_bank_port_1[0] && _zz_sram_2_banks_10_bank_port_2) begin
      sram_2_banks_10_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_10_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_10_bank_port_1[1] && _zz_sram_2_banks_10_bank_port_2) begin
      sram_2_banks_10_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_10_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_10_bank_port_1[2] && _zz_sram_2_banks_10_bank_port_2) begin
      sram_2_banks_10_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_10_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_10_bank_port_1[3] && _zz_sram_2_banks_10_bank_port_2) begin
      sram_2_banks_10_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_10_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_10_banksymbol_read <= sram_2_banks_10_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_10_banksymbol_read_1 <= sram_2_banks_10_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_10_banksymbol_read_2 <= sram_2_banks_10_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_10_banksymbol_read_3 <= sram_2_banks_10_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_11_bank_port1 = {_zz_sram_2_banks_11_banksymbol_read_3, _zz_sram_2_banks_11_banksymbol_read_2, _zz_sram_2_banks_11_banksymbol_read_1, _zz_sram_2_banks_11_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_2_banks_11_bank_port_1[0] && _zz_sram_2_banks_11_bank_port_2) begin
      sram_2_banks_11_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_11_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_11_bank_port_1[1] && _zz_sram_2_banks_11_bank_port_2) begin
      sram_2_banks_11_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_11_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_11_bank_port_1[2] && _zz_sram_2_banks_11_bank_port_2) begin
      sram_2_banks_11_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_11_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_11_bank_port_1[3] && _zz_sram_2_banks_11_bank_port_2) begin
      sram_2_banks_11_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_11_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_11_banksymbol_read <= sram_2_banks_11_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_11_banksymbol_read_1 <= sram_2_banks_11_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_11_banksymbol_read_2 <= sram_2_banks_11_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_11_banksymbol_read_3 <= sram_2_banks_11_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_12_bank_port1 = {_zz_sram_2_banks_12_banksymbol_read_3, _zz_sram_2_banks_12_banksymbol_read_2, _zz_sram_2_banks_12_banksymbol_read_1, _zz_sram_2_banks_12_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_2_banks_12_bank_port_1[0] && _zz_sram_2_banks_12_bank_port_2) begin
      sram_2_banks_12_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_12_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_12_bank_port_1[1] && _zz_sram_2_banks_12_bank_port_2) begin
      sram_2_banks_12_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_12_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_12_bank_port_1[2] && _zz_sram_2_banks_12_bank_port_2) begin
      sram_2_banks_12_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_12_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_12_bank_port_1[3] && _zz_sram_2_banks_12_bank_port_2) begin
      sram_2_banks_12_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_12_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_12_banksymbol_read <= sram_2_banks_12_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_12_banksymbol_read_1 <= sram_2_banks_12_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_12_banksymbol_read_2 <= sram_2_banks_12_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_12_banksymbol_read_3 <= sram_2_banks_12_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_13_bank_port1 = {_zz_sram_2_banks_13_banksymbol_read_3, _zz_sram_2_banks_13_banksymbol_read_2, _zz_sram_2_banks_13_banksymbol_read_1, _zz_sram_2_banks_13_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_2_banks_13_bank_port_1[0] && _zz_sram_2_banks_13_bank_port_2) begin
      sram_2_banks_13_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_13_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_13_bank_port_1[1] && _zz_sram_2_banks_13_bank_port_2) begin
      sram_2_banks_13_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_13_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_13_bank_port_1[2] && _zz_sram_2_banks_13_bank_port_2) begin
      sram_2_banks_13_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_13_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_13_bank_port_1[3] && _zz_sram_2_banks_13_bank_port_2) begin
      sram_2_banks_13_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_13_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_13_banksymbol_read <= sram_2_banks_13_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_13_banksymbol_read_1 <= sram_2_banks_13_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_13_banksymbol_read_2 <= sram_2_banks_13_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_13_banksymbol_read_3 <= sram_2_banks_13_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_14_bank_port1 = {_zz_sram_2_banks_14_banksymbol_read_3, _zz_sram_2_banks_14_banksymbol_read_2, _zz_sram_2_banks_14_banksymbol_read_1, _zz_sram_2_banks_14_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_2_banks_14_bank_port_1[0] && _zz_sram_2_banks_14_bank_port_2) begin
      sram_2_banks_14_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_14_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_14_bank_port_1[1] && _zz_sram_2_banks_14_bank_port_2) begin
      sram_2_banks_14_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_14_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_14_bank_port_1[2] && _zz_sram_2_banks_14_bank_port_2) begin
      sram_2_banks_14_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_14_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_14_bank_port_1[3] && _zz_sram_2_banks_14_bank_port_2) begin
      sram_2_banks_14_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_14_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_14_banksymbol_read <= sram_2_banks_14_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_14_banksymbol_read_1 <= sram_2_banks_14_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_14_banksymbol_read_2 <= sram_2_banks_14_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_14_banksymbol_read_3 <= sram_2_banks_14_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_2_banks_15_bank_port1 = {_zz_sram_2_banks_15_banksymbol_read_3, _zz_sram_2_banks_15_banksymbol_read_2, _zz_sram_2_banks_15_banksymbol_read_1, _zz_sram_2_banks_15_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_2_banks_15_bank_port_1[0] && _zz_sram_2_banks_15_bank_port_2) begin
      sram_2_banks_15_bank_symbol0[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_15_bank_port[7 : 0];
    end
    if(_zz_sram_2_banks_15_bank_port_1[1] && _zz_sram_2_banks_15_bank_port_2) begin
      sram_2_banks_15_bank_symbol1[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_15_bank_port[15 : 8];
    end
    if(_zz_sram_2_banks_15_bank_port_1[2] && _zz_sram_2_banks_15_bank_port_2) begin
      sram_2_banks_15_bank_symbol2[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_15_bank_port[23 : 16];
    end
    if(_zz_sram_2_banks_15_bank_port_1[3] && _zz_sram_2_banks_15_bank_port_2) begin
      sram_2_banks_15_bank_symbol3[sram_2_ports_cmd_payload_addr] <= _zz_sram_2_banks_15_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_2_ports_cmd_valid) begin
      _zz_sram_2_banks_15_banksymbol_read <= sram_2_banks_15_bank_symbol0[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_15_banksymbol_read_1 <= sram_2_banks_15_bank_symbol1[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_15_banksymbol_read_2 <= sram_2_banks_15_bank_symbol2[sram_2_ports_cmd_payload_addr];
      _zz_sram_2_banks_15_banksymbol_read_3 <= sram_2_banks_15_bank_symbol3[sram_2_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_0_bank_port1 = {_zz_sram_3_banks_0_banksymbol_read_3, _zz_sram_3_banks_0_banksymbol_read_2, _zz_sram_3_banks_0_banksymbol_read_1, _zz_sram_3_banks_0_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_3_banks_0_bank_port_1[0] && _zz_sram_3_banks_0_bank_port_2) begin
      sram_3_banks_0_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_0_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_0_bank_port_1[1] && _zz_sram_3_banks_0_bank_port_2) begin
      sram_3_banks_0_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_0_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_0_bank_port_1[2] && _zz_sram_3_banks_0_bank_port_2) begin
      sram_3_banks_0_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_0_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_0_bank_port_1[3] && _zz_sram_3_banks_0_bank_port_2) begin
      sram_3_banks_0_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_0_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_0_banksymbol_read <= sram_3_banks_0_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_0_banksymbol_read_1 <= sram_3_banks_0_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_0_banksymbol_read_2 <= sram_3_banks_0_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_0_banksymbol_read_3 <= sram_3_banks_0_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_1_bank_port1 = {_zz_sram_3_banks_1_banksymbol_read_3, _zz_sram_3_banks_1_banksymbol_read_2, _zz_sram_3_banks_1_banksymbol_read_1, _zz_sram_3_banks_1_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_3_banks_1_bank_port_1[0] && _zz_sram_3_banks_1_bank_port_2) begin
      sram_3_banks_1_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_1_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_1_bank_port_1[1] && _zz_sram_3_banks_1_bank_port_2) begin
      sram_3_banks_1_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_1_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_1_bank_port_1[2] && _zz_sram_3_banks_1_bank_port_2) begin
      sram_3_banks_1_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_1_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_1_bank_port_1[3] && _zz_sram_3_banks_1_bank_port_2) begin
      sram_3_banks_1_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_1_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_1_banksymbol_read <= sram_3_banks_1_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_1_banksymbol_read_1 <= sram_3_banks_1_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_1_banksymbol_read_2 <= sram_3_banks_1_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_1_banksymbol_read_3 <= sram_3_banks_1_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_2_bank_port1 = {_zz_sram_3_banks_2_banksymbol_read_3, _zz_sram_3_banks_2_banksymbol_read_2, _zz_sram_3_banks_2_banksymbol_read_1, _zz_sram_3_banks_2_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_3_banks_2_bank_port_1[0] && _zz_sram_3_banks_2_bank_port_2) begin
      sram_3_banks_2_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_2_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_2_bank_port_1[1] && _zz_sram_3_banks_2_bank_port_2) begin
      sram_3_banks_2_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_2_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_2_bank_port_1[2] && _zz_sram_3_banks_2_bank_port_2) begin
      sram_3_banks_2_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_2_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_2_bank_port_1[3] && _zz_sram_3_banks_2_bank_port_2) begin
      sram_3_banks_2_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_2_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_2_banksymbol_read <= sram_3_banks_2_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_2_banksymbol_read_1 <= sram_3_banks_2_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_2_banksymbol_read_2 <= sram_3_banks_2_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_2_banksymbol_read_3 <= sram_3_banks_2_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_3_bank_port1 = {_zz_sram_3_banks_3_banksymbol_read_3, _zz_sram_3_banks_3_banksymbol_read_2, _zz_sram_3_banks_3_banksymbol_read_1, _zz_sram_3_banks_3_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_3_banks_3_bank_port_1[0] && _zz_sram_3_banks_3_bank_port_2) begin
      sram_3_banks_3_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_3_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_3_bank_port_1[1] && _zz_sram_3_banks_3_bank_port_2) begin
      sram_3_banks_3_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_3_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_3_bank_port_1[2] && _zz_sram_3_banks_3_bank_port_2) begin
      sram_3_banks_3_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_3_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_3_bank_port_1[3] && _zz_sram_3_banks_3_bank_port_2) begin
      sram_3_banks_3_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_3_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_3_banksymbol_read <= sram_3_banks_3_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_3_banksymbol_read_1 <= sram_3_banks_3_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_3_banksymbol_read_2 <= sram_3_banks_3_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_3_banksymbol_read_3 <= sram_3_banks_3_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_4_bank_port1 = {_zz_sram_3_banks_4_banksymbol_read_3, _zz_sram_3_banks_4_banksymbol_read_2, _zz_sram_3_banks_4_banksymbol_read_1, _zz_sram_3_banks_4_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_3_banks_4_bank_port_1[0] && _zz_sram_3_banks_4_bank_port_2) begin
      sram_3_banks_4_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_4_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_4_bank_port_1[1] && _zz_sram_3_banks_4_bank_port_2) begin
      sram_3_banks_4_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_4_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_4_bank_port_1[2] && _zz_sram_3_banks_4_bank_port_2) begin
      sram_3_banks_4_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_4_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_4_bank_port_1[3] && _zz_sram_3_banks_4_bank_port_2) begin
      sram_3_banks_4_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_4_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_4_banksymbol_read <= sram_3_banks_4_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_4_banksymbol_read_1 <= sram_3_banks_4_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_4_banksymbol_read_2 <= sram_3_banks_4_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_4_banksymbol_read_3 <= sram_3_banks_4_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_5_bank_port1 = {_zz_sram_3_banks_5_banksymbol_read_3, _zz_sram_3_banks_5_banksymbol_read_2, _zz_sram_3_banks_5_banksymbol_read_1, _zz_sram_3_banks_5_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_3_banks_5_bank_port_1[0] && _zz_sram_3_banks_5_bank_port_2) begin
      sram_3_banks_5_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_5_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_5_bank_port_1[1] && _zz_sram_3_banks_5_bank_port_2) begin
      sram_3_banks_5_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_5_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_5_bank_port_1[2] && _zz_sram_3_banks_5_bank_port_2) begin
      sram_3_banks_5_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_5_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_5_bank_port_1[3] && _zz_sram_3_banks_5_bank_port_2) begin
      sram_3_banks_5_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_5_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_5_banksymbol_read <= sram_3_banks_5_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_5_banksymbol_read_1 <= sram_3_banks_5_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_5_banksymbol_read_2 <= sram_3_banks_5_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_5_banksymbol_read_3 <= sram_3_banks_5_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_6_bank_port1 = {_zz_sram_3_banks_6_banksymbol_read_3, _zz_sram_3_banks_6_banksymbol_read_2, _zz_sram_3_banks_6_banksymbol_read_1, _zz_sram_3_banks_6_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_3_banks_6_bank_port_1[0] && _zz_sram_3_banks_6_bank_port_2) begin
      sram_3_banks_6_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_6_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_6_bank_port_1[1] && _zz_sram_3_banks_6_bank_port_2) begin
      sram_3_banks_6_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_6_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_6_bank_port_1[2] && _zz_sram_3_banks_6_bank_port_2) begin
      sram_3_banks_6_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_6_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_6_bank_port_1[3] && _zz_sram_3_banks_6_bank_port_2) begin
      sram_3_banks_6_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_6_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_6_banksymbol_read <= sram_3_banks_6_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_6_banksymbol_read_1 <= sram_3_banks_6_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_6_banksymbol_read_2 <= sram_3_banks_6_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_6_banksymbol_read_3 <= sram_3_banks_6_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_7_bank_port1 = {_zz_sram_3_banks_7_banksymbol_read_3, _zz_sram_3_banks_7_banksymbol_read_2, _zz_sram_3_banks_7_banksymbol_read_1, _zz_sram_3_banks_7_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_3_banks_7_bank_port_1[0] && _zz_sram_3_banks_7_bank_port_2) begin
      sram_3_banks_7_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_7_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_7_bank_port_1[1] && _zz_sram_3_banks_7_bank_port_2) begin
      sram_3_banks_7_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_7_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_7_bank_port_1[2] && _zz_sram_3_banks_7_bank_port_2) begin
      sram_3_banks_7_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_7_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_7_bank_port_1[3] && _zz_sram_3_banks_7_bank_port_2) begin
      sram_3_banks_7_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_7_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_7_banksymbol_read <= sram_3_banks_7_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_7_banksymbol_read_1 <= sram_3_banks_7_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_7_banksymbol_read_2 <= sram_3_banks_7_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_7_banksymbol_read_3 <= sram_3_banks_7_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_8_bank_port1 = {_zz_sram_3_banks_8_banksymbol_read_3, _zz_sram_3_banks_8_banksymbol_read_2, _zz_sram_3_banks_8_banksymbol_read_1, _zz_sram_3_banks_8_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_3_banks_8_bank_port_1[0] && _zz_sram_3_banks_8_bank_port_2) begin
      sram_3_banks_8_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_8_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_8_bank_port_1[1] && _zz_sram_3_banks_8_bank_port_2) begin
      sram_3_banks_8_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_8_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_8_bank_port_1[2] && _zz_sram_3_banks_8_bank_port_2) begin
      sram_3_banks_8_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_8_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_8_bank_port_1[3] && _zz_sram_3_banks_8_bank_port_2) begin
      sram_3_banks_8_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_8_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_8_banksymbol_read <= sram_3_banks_8_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_8_banksymbol_read_1 <= sram_3_banks_8_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_8_banksymbol_read_2 <= sram_3_banks_8_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_8_banksymbol_read_3 <= sram_3_banks_8_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_9_bank_port1 = {_zz_sram_3_banks_9_banksymbol_read_3, _zz_sram_3_banks_9_banksymbol_read_2, _zz_sram_3_banks_9_banksymbol_read_1, _zz_sram_3_banks_9_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_3_banks_9_bank_port_1[0] && _zz_sram_3_banks_9_bank_port_2) begin
      sram_3_banks_9_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_9_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_9_bank_port_1[1] && _zz_sram_3_banks_9_bank_port_2) begin
      sram_3_banks_9_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_9_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_9_bank_port_1[2] && _zz_sram_3_banks_9_bank_port_2) begin
      sram_3_banks_9_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_9_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_9_bank_port_1[3] && _zz_sram_3_banks_9_bank_port_2) begin
      sram_3_banks_9_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_9_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_9_banksymbol_read <= sram_3_banks_9_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_9_banksymbol_read_1 <= sram_3_banks_9_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_9_banksymbol_read_2 <= sram_3_banks_9_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_9_banksymbol_read_3 <= sram_3_banks_9_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_10_bank_port1 = {_zz_sram_3_banks_10_banksymbol_read_3, _zz_sram_3_banks_10_banksymbol_read_2, _zz_sram_3_banks_10_banksymbol_read_1, _zz_sram_3_banks_10_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_3_banks_10_bank_port_1[0] && _zz_sram_3_banks_10_bank_port_2) begin
      sram_3_banks_10_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_10_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_10_bank_port_1[1] && _zz_sram_3_banks_10_bank_port_2) begin
      sram_3_banks_10_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_10_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_10_bank_port_1[2] && _zz_sram_3_banks_10_bank_port_2) begin
      sram_3_banks_10_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_10_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_10_bank_port_1[3] && _zz_sram_3_banks_10_bank_port_2) begin
      sram_3_banks_10_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_10_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_10_banksymbol_read <= sram_3_banks_10_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_10_banksymbol_read_1 <= sram_3_banks_10_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_10_banksymbol_read_2 <= sram_3_banks_10_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_10_banksymbol_read_3 <= sram_3_banks_10_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_11_bank_port1 = {_zz_sram_3_banks_11_banksymbol_read_3, _zz_sram_3_banks_11_banksymbol_read_2, _zz_sram_3_banks_11_banksymbol_read_1, _zz_sram_3_banks_11_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_3_banks_11_bank_port_1[0] && _zz_sram_3_banks_11_bank_port_2) begin
      sram_3_banks_11_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_11_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_11_bank_port_1[1] && _zz_sram_3_banks_11_bank_port_2) begin
      sram_3_banks_11_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_11_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_11_bank_port_1[2] && _zz_sram_3_banks_11_bank_port_2) begin
      sram_3_banks_11_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_11_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_11_bank_port_1[3] && _zz_sram_3_banks_11_bank_port_2) begin
      sram_3_banks_11_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_11_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_11_banksymbol_read <= sram_3_banks_11_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_11_banksymbol_read_1 <= sram_3_banks_11_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_11_banksymbol_read_2 <= sram_3_banks_11_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_11_banksymbol_read_3 <= sram_3_banks_11_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_12_bank_port1 = {_zz_sram_3_banks_12_banksymbol_read_3, _zz_sram_3_banks_12_banksymbol_read_2, _zz_sram_3_banks_12_banksymbol_read_1, _zz_sram_3_banks_12_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_3_banks_12_bank_port_1[0] && _zz_sram_3_banks_12_bank_port_2) begin
      sram_3_banks_12_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_12_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_12_bank_port_1[1] && _zz_sram_3_banks_12_bank_port_2) begin
      sram_3_banks_12_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_12_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_12_bank_port_1[2] && _zz_sram_3_banks_12_bank_port_2) begin
      sram_3_banks_12_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_12_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_12_bank_port_1[3] && _zz_sram_3_banks_12_bank_port_2) begin
      sram_3_banks_12_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_12_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_12_banksymbol_read <= sram_3_banks_12_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_12_banksymbol_read_1 <= sram_3_banks_12_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_12_banksymbol_read_2 <= sram_3_banks_12_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_12_banksymbol_read_3 <= sram_3_banks_12_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_13_bank_port1 = {_zz_sram_3_banks_13_banksymbol_read_3, _zz_sram_3_banks_13_banksymbol_read_2, _zz_sram_3_banks_13_banksymbol_read_1, _zz_sram_3_banks_13_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_3_banks_13_bank_port_1[0] && _zz_sram_3_banks_13_bank_port_2) begin
      sram_3_banks_13_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_13_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_13_bank_port_1[1] && _zz_sram_3_banks_13_bank_port_2) begin
      sram_3_banks_13_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_13_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_13_bank_port_1[2] && _zz_sram_3_banks_13_bank_port_2) begin
      sram_3_banks_13_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_13_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_13_bank_port_1[3] && _zz_sram_3_banks_13_bank_port_2) begin
      sram_3_banks_13_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_13_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_13_banksymbol_read <= sram_3_banks_13_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_13_banksymbol_read_1 <= sram_3_banks_13_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_13_banksymbol_read_2 <= sram_3_banks_13_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_13_banksymbol_read_3 <= sram_3_banks_13_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_14_bank_port1 = {_zz_sram_3_banks_14_banksymbol_read_3, _zz_sram_3_banks_14_banksymbol_read_2, _zz_sram_3_banks_14_banksymbol_read_1, _zz_sram_3_banks_14_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_3_banks_14_bank_port_1[0] && _zz_sram_3_banks_14_bank_port_2) begin
      sram_3_banks_14_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_14_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_14_bank_port_1[1] && _zz_sram_3_banks_14_bank_port_2) begin
      sram_3_banks_14_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_14_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_14_bank_port_1[2] && _zz_sram_3_banks_14_bank_port_2) begin
      sram_3_banks_14_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_14_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_14_bank_port_1[3] && _zz_sram_3_banks_14_bank_port_2) begin
      sram_3_banks_14_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_14_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_14_banksymbol_read <= sram_3_banks_14_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_14_banksymbol_read_1 <= sram_3_banks_14_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_14_banksymbol_read_2 <= sram_3_banks_14_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_14_banksymbol_read_3 <= sram_3_banks_14_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    _zz_sram_3_banks_15_bank_port1 = {_zz_sram_3_banks_15_banksymbol_read_3, _zz_sram_3_banks_15_banksymbol_read_2, _zz_sram_3_banks_15_banksymbol_read_1, _zz_sram_3_banks_15_banksymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_sram_3_banks_15_bank_port_1[0] && _zz_sram_3_banks_15_bank_port_2) begin
      sram_3_banks_15_bank_symbol0[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_15_bank_port[7 : 0];
    end
    if(_zz_sram_3_banks_15_bank_port_1[1] && _zz_sram_3_banks_15_bank_port_2) begin
      sram_3_banks_15_bank_symbol1[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_15_bank_port[15 : 8];
    end
    if(_zz_sram_3_banks_15_bank_port_1[2] && _zz_sram_3_banks_15_bank_port_2) begin
      sram_3_banks_15_bank_symbol2[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_15_bank_port[23 : 16];
    end
    if(_zz_sram_3_banks_15_bank_port_1[3] && _zz_sram_3_banks_15_bank_port_2) begin
      sram_3_banks_15_bank_symbol3[sram_3_ports_cmd_payload_addr] <= _zz_sram_3_banks_15_bank_port[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(sram_3_ports_cmd_valid) begin
      _zz_sram_3_banks_15_banksymbol_read <= sram_3_banks_15_bank_symbol0[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_15_banksymbol_read_1 <= sram_3_banks_15_bank_symbol1[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_15_banksymbol_read_2 <= sram_3_banks_15_bank_symbol2[sram_3_ports_cmd_payload_addr];
      _zz_sram_3_banks_15_banksymbol_read_3 <= sram_3_banks_15_bank_symbol3[sram_3_ports_cmd_payload_addr];
    end
  end

  always @(*) begin
    sram_0_ports_rsp_payload_data[31 : 0] = _zz_sram_0_banks_0_bank_port1;
    sram_0_ports_rsp_payload_data[63 : 32] = _zz_sram_0_banks_1_bank_port1;
    sram_0_ports_rsp_payload_data[95 : 64] = _zz_sram_0_banks_2_bank_port1;
    sram_0_ports_rsp_payload_data[127 : 96] = _zz_sram_0_banks_3_bank_port1;
    sram_0_ports_rsp_payload_data[159 : 128] = _zz_sram_0_banks_4_bank_port1;
    sram_0_ports_rsp_payload_data[191 : 160] = _zz_sram_0_banks_5_bank_port1;
    sram_0_ports_rsp_payload_data[223 : 192] = _zz_sram_0_banks_6_bank_port1;
    sram_0_ports_rsp_payload_data[255 : 224] = _zz_sram_0_banks_7_bank_port1;
    sram_0_ports_rsp_payload_data[287 : 256] = _zz_sram_0_banks_8_bank_port1;
    sram_0_ports_rsp_payload_data[319 : 288] = _zz_sram_0_banks_9_bank_port1;
    sram_0_ports_rsp_payload_data[351 : 320] = _zz_sram_0_banks_10_bank_port1;
    sram_0_ports_rsp_payload_data[383 : 352] = _zz_sram_0_banks_11_bank_port1;
    sram_0_ports_rsp_payload_data[415 : 384] = _zz_sram_0_banks_12_bank_port1;
    sram_0_ports_rsp_payload_data[447 : 416] = _zz_sram_0_banks_13_bank_port1;
    sram_0_ports_rsp_payload_data[479 : 448] = _zz_sram_0_banks_14_bank_port1;
    sram_0_ports_rsp_payload_data[511 : 480] = _zz_sram_0_banks_15_bank_port1;
  end

  assign when_SramBanks_l66 = (sram_0_ports_cmd_valid && (sram_0_ports_cmd_payload_wen == 16'h0));
  assign sram_0_ports_rsp_valid = _zz_sram_0_ports_rsp_valid;
  always @(*) begin
    sram_1_ports_rsp_payload_data[31 : 0] = _zz_sram_1_banks_0_bank_port1;
    sram_1_ports_rsp_payload_data[63 : 32] = _zz_sram_1_banks_1_bank_port1;
    sram_1_ports_rsp_payload_data[95 : 64] = _zz_sram_1_banks_2_bank_port1;
    sram_1_ports_rsp_payload_data[127 : 96] = _zz_sram_1_banks_3_bank_port1;
    sram_1_ports_rsp_payload_data[159 : 128] = _zz_sram_1_banks_4_bank_port1;
    sram_1_ports_rsp_payload_data[191 : 160] = _zz_sram_1_banks_5_bank_port1;
    sram_1_ports_rsp_payload_data[223 : 192] = _zz_sram_1_banks_6_bank_port1;
    sram_1_ports_rsp_payload_data[255 : 224] = _zz_sram_1_banks_7_bank_port1;
    sram_1_ports_rsp_payload_data[287 : 256] = _zz_sram_1_banks_8_bank_port1;
    sram_1_ports_rsp_payload_data[319 : 288] = _zz_sram_1_banks_9_bank_port1;
    sram_1_ports_rsp_payload_data[351 : 320] = _zz_sram_1_banks_10_bank_port1;
    sram_1_ports_rsp_payload_data[383 : 352] = _zz_sram_1_banks_11_bank_port1;
    sram_1_ports_rsp_payload_data[415 : 384] = _zz_sram_1_banks_12_bank_port1;
    sram_1_ports_rsp_payload_data[447 : 416] = _zz_sram_1_banks_13_bank_port1;
    sram_1_ports_rsp_payload_data[479 : 448] = _zz_sram_1_banks_14_bank_port1;
    sram_1_ports_rsp_payload_data[511 : 480] = _zz_sram_1_banks_15_bank_port1;
  end

  assign when_SramBanks_l66_1 = (sram_1_ports_cmd_valid && (sram_1_ports_cmd_payload_wen == 16'h0));
  assign sram_1_ports_rsp_valid = _zz_sram_1_ports_rsp_valid;
  always @(*) begin
    sram_2_ports_rsp_payload_data[31 : 0] = _zz_sram_2_banks_0_bank_port1;
    sram_2_ports_rsp_payload_data[63 : 32] = _zz_sram_2_banks_1_bank_port1;
    sram_2_ports_rsp_payload_data[95 : 64] = _zz_sram_2_banks_2_bank_port1;
    sram_2_ports_rsp_payload_data[127 : 96] = _zz_sram_2_banks_3_bank_port1;
    sram_2_ports_rsp_payload_data[159 : 128] = _zz_sram_2_banks_4_bank_port1;
    sram_2_ports_rsp_payload_data[191 : 160] = _zz_sram_2_banks_5_bank_port1;
    sram_2_ports_rsp_payload_data[223 : 192] = _zz_sram_2_banks_6_bank_port1;
    sram_2_ports_rsp_payload_data[255 : 224] = _zz_sram_2_banks_7_bank_port1;
    sram_2_ports_rsp_payload_data[287 : 256] = _zz_sram_2_banks_8_bank_port1;
    sram_2_ports_rsp_payload_data[319 : 288] = _zz_sram_2_banks_9_bank_port1;
    sram_2_ports_rsp_payload_data[351 : 320] = _zz_sram_2_banks_10_bank_port1;
    sram_2_ports_rsp_payload_data[383 : 352] = _zz_sram_2_banks_11_bank_port1;
    sram_2_ports_rsp_payload_data[415 : 384] = _zz_sram_2_banks_12_bank_port1;
    sram_2_ports_rsp_payload_data[447 : 416] = _zz_sram_2_banks_13_bank_port1;
    sram_2_ports_rsp_payload_data[479 : 448] = _zz_sram_2_banks_14_bank_port1;
    sram_2_ports_rsp_payload_data[511 : 480] = _zz_sram_2_banks_15_bank_port1;
  end

  assign when_SramBanks_l66_2 = (sram_2_ports_cmd_valid && (sram_2_ports_cmd_payload_wen == 16'h0));
  assign sram_2_ports_rsp_valid = _zz_sram_2_ports_rsp_valid;
  always @(*) begin
    sram_3_ports_rsp_payload_data[31 : 0] = _zz_sram_3_banks_0_bank_port1;
    sram_3_ports_rsp_payload_data[63 : 32] = _zz_sram_3_banks_1_bank_port1;
    sram_3_ports_rsp_payload_data[95 : 64] = _zz_sram_3_banks_2_bank_port1;
    sram_3_ports_rsp_payload_data[127 : 96] = _zz_sram_3_banks_3_bank_port1;
    sram_3_ports_rsp_payload_data[159 : 128] = _zz_sram_3_banks_4_bank_port1;
    sram_3_ports_rsp_payload_data[191 : 160] = _zz_sram_3_banks_5_bank_port1;
    sram_3_ports_rsp_payload_data[223 : 192] = _zz_sram_3_banks_6_bank_port1;
    sram_3_ports_rsp_payload_data[255 : 224] = _zz_sram_3_banks_7_bank_port1;
    sram_3_ports_rsp_payload_data[287 : 256] = _zz_sram_3_banks_8_bank_port1;
    sram_3_ports_rsp_payload_data[319 : 288] = _zz_sram_3_banks_9_bank_port1;
    sram_3_ports_rsp_payload_data[351 : 320] = _zz_sram_3_banks_10_bank_port1;
    sram_3_ports_rsp_payload_data[383 : 352] = _zz_sram_3_banks_11_bank_port1;
    sram_3_ports_rsp_payload_data[415 : 384] = _zz_sram_3_banks_12_bank_port1;
    sram_3_ports_rsp_payload_data[447 : 416] = _zz_sram_3_banks_13_bank_port1;
    sram_3_ports_rsp_payload_data[479 : 448] = _zz_sram_3_banks_14_bank_port1;
    sram_3_ports_rsp_payload_data[511 : 480] = _zz_sram_3_banks_15_bank_port1;
  end

  assign when_SramBanks_l66_3 = (sram_3_ports_cmd_valid && (sram_3_ports_cmd_payload_wen == 16'h0));
  assign sram_3_ports_rsp_valid = _zz_sram_3_ports_rsp_valid;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _zz_sram_0_ports_rsp_valid <= 1'b0;
      _zz_sram_1_ports_rsp_valid <= 1'b0;
      _zz_sram_2_ports_rsp_valid <= 1'b0;
      _zz_sram_3_ports_rsp_valid <= 1'b0;
    end else begin
      if(when_SramBanks_l66) begin
        _zz_sram_0_ports_rsp_valid <= 1'b1;
      end else begin
        _zz_sram_0_ports_rsp_valid <= 1'b0;
      end
      if(when_SramBanks_l66_1) begin
        _zz_sram_1_ports_rsp_valid <= 1'b1;
      end else begin
        _zz_sram_1_ports_rsp_valid <= 1'b0;
      end
      if(when_SramBanks_l66_2) begin
        _zz_sram_2_ports_rsp_valid <= 1'b1;
      end else begin
        _zz_sram_2_ports_rsp_valid <= 1'b0;
      end
      if(when_SramBanks_l66_3) begin
        _zz_sram_3_ports_rsp_valid <= 1'b1;
      end else begin
        _zz_sram_3_ports_rsp_valid <= 1'b0;
      end
    end
  end


endmodule

module ICache (
  input               flush,
  input               cpu_cmd_valid,
  output              cpu_cmd_ready,
  input      [63:0]   cpu_cmd_payload_addr,
  output              cpu_rsp_valid,
  output     [31:0]   cpu_rsp_payload_data,
  output reg          sram_0_ports_cmd_valid,
  output reg [6:0]    sram_0_ports_cmd_payload_addr,
  output reg [15:0]   sram_0_ports_cmd_payload_wen,
  output reg [511:0]  sram_0_ports_cmd_payload_wdata,
  output reg [63:0]   sram_0_ports_cmd_payload_wstrb,
  input               sram_0_ports_rsp_valid,
  input      [511:0]  sram_0_ports_rsp_payload_data,
  output reg          sram_1_ports_cmd_valid,
  output reg [6:0]    sram_1_ports_cmd_payload_addr,
  output reg [15:0]   sram_1_ports_cmd_payload_wen,
  output reg [511:0]  sram_1_ports_cmd_payload_wdata,
  output reg [63:0]   sram_1_ports_cmd_payload_wstrb,
  input               sram_1_ports_rsp_valid,
  input      [511:0]  sram_1_ports_rsp_payload_data,
  output reg          sram_2_ports_cmd_valid,
  output reg [6:0]    sram_2_ports_cmd_payload_addr,
  output reg [15:0]   sram_2_ports_cmd_payload_wen,
  output reg [511:0]  sram_2_ports_cmd_payload_wdata,
  output reg [63:0]   sram_2_ports_cmd_payload_wstrb,
  input               sram_2_ports_rsp_valid,
  input      [511:0]  sram_2_ports_rsp_payload_data,
  output reg          sram_3_ports_cmd_valid,
  output reg [6:0]    sram_3_ports_cmd_payload_addr,
  output reg [15:0]   sram_3_ports_cmd_payload_wen,
  output reg [511:0]  sram_3_ports_cmd_payload_wdata,
  output reg [63:0]   sram_3_ports_cmd_payload_wstrb,
  input               sram_3_ports_rsp_valid,
  input      [511:0]  sram_3_ports_rsp_payload_data,
  output              sram_4_ports_cmd_valid,
  output     [6:0]    sram_4_ports_cmd_payload_addr,
  output     [15:0]   sram_4_ports_cmd_payload_wen,
  output     [511:0]  sram_4_ports_cmd_payload_wdata,
  output     [63:0]   sram_4_ports_cmd_payload_wstrb,
  input               sram_4_ports_rsp_valid,
  input      [511:0]  sram_4_ports_rsp_payload_data,
  output              sram_5_ports_cmd_valid,
  output     [6:0]    sram_5_ports_cmd_payload_addr,
  output     [15:0]   sram_5_ports_cmd_payload_wen,
  output     [511:0]  sram_5_ports_cmd_payload_wdata,
  output     [63:0]   sram_5_ports_cmd_payload_wstrb,
  input               sram_5_ports_rsp_valid,
  input      [511:0]  sram_5_ports_rsp_payload_data,
  output              sram_6_ports_cmd_valid,
  output     [6:0]    sram_6_ports_cmd_payload_addr,
  output     [15:0]   sram_6_ports_cmd_payload_wen,
  output     [511:0]  sram_6_ports_cmd_payload_wdata,
  output     [63:0]   sram_6_ports_cmd_payload_wstrb,
  input               sram_6_ports_rsp_valid,
  input      [511:0]  sram_6_ports_rsp_payload_data,
  output              sram_7_ports_cmd_valid,
  output     [6:0]    sram_7_ports_cmd_payload_addr,
  output     [15:0]   sram_7_ports_cmd_payload_wen,
  output     [511:0]  sram_7_ports_cmd_payload_wdata,
  output     [63:0]   sram_7_ports_cmd_payload_wstrb,
  input               sram_7_ports_rsp_valid,
  input      [511:0]  sram_7_ports_rsp_payload_data,
  output              sram_8_ports_cmd_valid,
  output     [6:0]    sram_8_ports_cmd_payload_addr,
  output     [15:0]   sram_8_ports_cmd_payload_wen,
  output     [511:0]  sram_8_ports_cmd_payload_wdata,
  output     [63:0]   sram_8_ports_cmd_payload_wstrb,
  input               sram_8_ports_rsp_valid,
  input      [511:0]  sram_8_ports_rsp_payload_data,
  output              sram_9_ports_cmd_valid,
  output     [6:0]    sram_9_ports_cmd_payload_addr,
  output     [15:0]   sram_9_ports_cmd_payload_wen,
  output     [511:0]  sram_9_ports_cmd_payload_wdata,
  output     [63:0]   sram_9_ports_cmd_payload_wstrb,
  input               sram_9_ports_rsp_valid,
  input      [511:0]  sram_9_ports_rsp_payload_data,
  output              sram_10_ports_cmd_valid,
  output     [6:0]    sram_10_ports_cmd_payload_addr,
  output     [15:0]   sram_10_ports_cmd_payload_wen,
  output     [511:0]  sram_10_ports_cmd_payload_wdata,
  output     [63:0]   sram_10_ports_cmd_payload_wstrb,
  input               sram_10_ports_rsp_valid,
  input      [511:0]  sram_10_ports_rsp_payload_data,
  output              sram_11_ports_cmd_valid,
  output     [6:0]    sram_11_ports_cmd_payload_addr,
  output     [15:0]   sram_11_ports_cmd_payload_wen,
  output     [511:0]  sram_11_ports_cmd_payload_wdata,
  output     [63:0]   sram_11_ports_cmd_payload_wstrb,
  input               sram_11_ports_rsp_valid,
  input      [511:0]  sram_11_ports_rsp_payload_data,
  output              sram_12_ports_cmd_valid,
  output     [6:0]    sram_12_ports_cmd_payload_addr,
  output     [15:0]   sram_12_ports_cmd_payload_wen,
  output     [511:0]  sram_12_ports_cmd_payload_wdata,
  output     [63:0]   sram_12_ports_cmd_payload_wstrb,
  input               sram_12_ports_rsp_valid,
  input      [511:0]  sram_12_ports_rsp_payload_data,
  output              sram_13_ports_cmd_valid,
  output     [6:0]    sram_13_ports_cmd_payload_addr,
  output     [15:0]   sram_13_ports_cmd_payload_wen,
  output     [511:0]  sram_13_ports_cmd_payload_wdata,
  output     [63:0]   sram_13_ports_cmd_payload_wstrb,
  input               sram_13_ports_rsp_valid,
  input      [511:0]  sram_13_ports_rsp_payload_data,
  output              sram_14_ports_cmd_valid,
  output     [6:0]    sram_14_ports_cmd_payload_addr,
  output     [15:0]   sram_14_ports_cmd_payload_wen,
  output     [511:0]  sram_14_ports_cmd_payload_wdata,
  output     [63:0]   sram_14_ports_cmd_payload_wstrb,
  input               sram_14_ports_rsp_valid,
  input      [511:0]  sram_14_ports_rsp_payload_data,
  output              sram_15_ports_cmd_valid,
  output     [6:0]    sram_15_ports_cmd_payload_addr,
  output     [15:0]   sram_15_ports_cmd_payload_wen,
  output     [511:0]  sram_15_ports_cmd_payload_wdata,
  output     [63:0]   sram_15_ports_cmd_payload_wstrb,
  input               sram_15_ports_rsp_valid,
  input      [511:0]  sram_15_ports_rsp_payload_data,
  output              next_level_cmd_valid,
  input               next_level_cmd_ready,
  output     [63:0]   next_level_cmd_payload_addr,
  output     [3:0]    next_level_cmd_payload_len,
  output     [2:0]    next_level_cmd_payload_size,
  input               next_level_rsp_valid,
  input      [63:0]   next_level_rsp_payload_data,
  input               clk,
  input               reset
);

  wire       [6:0]    _zz_flush_cnt_valueNext;
  wire       [0:0]    _zz_flush_cnt_valueNext_1;
  wire       [2:0]    _zz_next_level_data_cnt_valueNext;
  wire       [0:0]    _zz_next_level_data_cnt_valueNext_1;
  wire       [7:0]    _zz__zz_cache_hit_gnt_0_3;
  wire       [7:0]    _zz__zz_cache_hit_gnt_0_3_1;
  wire       [3:0]    _zz__zz_cache_hit_gnt_0_3_2;
  wire       [7:0]    _zz__zz_cache_invld_gnt_0_3;
  wire       [7:0]    _zz__zz_cache_invld_gnt_0_3_1;
  wire       [3:0]    _zz__zz_cache_invld_gnt_0_3_2;
  wire       [7:0]    _zz__zz_cache_victim_gnt_0_3;
  wire       [7:0]    _zz__zz_cache_victim_gnt_0_3_1;
  wire       [3:0]    _zz__zz_cache_victim_gnt_0_3_2;
  reg        [50:0]   _zz_cache_tag_0;
  reg                 _zz_cache_hit_0;
  reg                 _zz_cache_mru_0;
  reg                 _zz_cache_invld_d1_0;
  reg                 _zz_cache_lru_d1_0;
  wire       [4:0]    _zz_sram_0_ports_cmd_payload_wen_1;
  wire       [9:0]    _zz_sram_0_ports_cmd_payload_wdata;
  wire       [9:0]    _zz_sram_0_ports_cmd_payload_wstrb;
  wire       [9:0]    _zz_sram_0_ports_cmd_payload_wstrb_1;
  reg        [50:0]   _zz_cache_tag_1;
  reg                 _zz_cache_hit_1;
  reg                 _zz_cache_mru_1;
  reg                 _zz_cache_invld_d1_1;
  reg                 _zz_cache_lru_d1_1;
  wire       [4:0]    _zz_sram_1_ports_cmd_payload_wen_1;
  wire       [9:0]    _zz_sram_1_ports_cmd_payload_wdata;
  wire       [9:0]    _zz_sram_1_ports_cmd_payload_wstrb;
  wire       [9:0]    _zz_sram_1_ports_cmd_payload_wstrb_1;
  reg        [50:0]   _zz_cache_tag_2;
  reg                 _zz_cache_hit_2;
  reg                 _zz_cache_mru_2;
  reg                 _zz_cache_invld_d1_2;
  reg                 _zz_cache_lru_d1_2;
  wire       [4:0]    _zz_sram_2_ports_cmd_payload_wen_1;
  wire       [9:0]    _zz_sram_2_ports_cmd_payload_wdata;
  wire       [9:0]    _zz_sram_2_ports_cmd_payload_wstrb;
  wire       [9:0]    _zz_sram_2_ports_cmd_payload_wstrb_1;
  reg        [50:0]   _zz_cache_tag_3;
  reg                 _zz_cache_hit_3;
  reg                 _zz_cache_mru_3;
  reg                 _zz_cache_invld_d1_3;
  reg                 _zz_cache_lru_d1_3;
  wire       [4:0]    _zz_sram_3_ports_cmd_payload_wen_1;
  wire       [9:0]    _zz_sram_3_ports_cmd_payload_wdata;
  wire       [9:0]    _zz_sram_3_ports_cmd_payload_wstrb;
  wire       [9:0]    _zz_sram_3_ports_cmd_payload_wstrb_1;
  reg        [511:0]  _zz__zz_cpu_rsp_payload_data;
  reg        [511:0]  _zz__zz_cpu_rsp_payload_data_1;
  reg        [31:0]   _zz_cpu_rsp_payload_data_2;
  reg        [31:0]   _zz_cpu_rsp_payload_data_3;
  reg                 _zz_cpu_rsp_valid;
  reg                 _zz_cpu_rsp_valid_1;
  reg                 ways_0_metas_0_vld;
  reg        [50:0]   ways_0_metas_0_tag;
  reg                 ways_0_metas_0_mru;
  reg                 ways_0_metas_1_vld;
  reg        [50:0]   ways_0_metas_1_tag;
  reg                 ways_0_metas_1_mru;
  reg                 ways_0_metas_2_vld;
  reg        [50:0]   ways_0_metas_2_tag;
  reg                 ways_0_metas_2_mru;
  reg                 ways_0_metas_3_vld;
  reg        [50:0]   ways_0_metas_3_tag;
  reg                 ways_0_metas_3_mru;
  reg                 ways_0_metas_4_vld;
  reg        [50:0]   ways_0_metas_4_tag;
  reg                 ways_0_metas_4_mru;
  reg                 ways_0_metas_5_vld;
  reg        [50:0]   ways_0_metas_5_tag;
  reg                 ways_0_metas_5_mru;
  reg                 ways_0_metas_6_vld;
  reg        [50:0]   ways_0_metas_6_tag;
  reg                 ways_0_metas_6_mru;
  reg                 ways_0_metas_7_vld;
  reg        [50:0]   ways_0_metas_7_tag;
  reg                 ways_0_metas_7_mru;
  reg                 ways_0_metas_8_vld;
  reg        [50:0]   ways_0_metas_8_tag;
  reg                 ways_0_metas_8_mru;
  reg                 ways_0_metas_9_vld;
  reg        [50:0]   ways_0_metas_9_tag;
  reg                 ways_0_metas_9_mru;
  reg                 ways_0_metas_10_vld;
  reg        [50:0]   ways_0_metas_10_tag;
  reg                 ways_0_metas_10_mru;
  reg                 ways_0_metas_11_vld;
  reg        [50:0]   ways_0_metas_11_tag;
  reg                 ways_0_metas_11_mru;
  reg                 ways_0_metas_12_vld;
  reg        [50:0]   ways_0_metas_12_tag;
  reg                 ways_0_metas_12_mru;
  reg                 ways_0_metas_13_vld;
  reg        [50:0]   ways_0_metas_13_tag;
  reg                 ways_0_metas_13_mru;
  reg                 ways_0_metas_14_vld;
  reg        [50:0]   ways_0_metas_14_tag;
  reg                 ways_0_metas_14_mru;
  reg                 ways_0_metas_15_vld;
  reg        [50:0]   ways_0_metas_15_tag;
  reg                 ways_0_metas_15_mru;
  reg                 ways_0_metas_16_vld;
  reg        [50:0]   ways_0_metas_16_tag;
  reg                 ways_0_metas_16_mru;
  reg                 ways_0_metas_17_vld;
  reg        [50:0]   ways_0_metas_17_tag;
  reg                 ways_0_metas_17_mru;
  reg                 ways_0_metas_18_vld;
  reg        [50:0]   ways_0_metas_18_tag;
  reg                 ways_0_metas_18_mru;
  reg                 ways_0_metas_19_vld;
  reg        [50:0]   ways_0_metas_19_tag;
  reg                 ways_0_metas_19_mru;
  reg                 ways_0_metas_20_vld;
  reg        [50:0]   ways_0_metas_20_tag;
  reg                 ways_0_metas_20_mru;
  reg                 ways_0_metas_21_vld;
  reg        [50:0]   ways_0_metas_21_tag;
  reg                 ways_0_metas_21_mru;
  reg                 ways_0_metas_22_vld;
  reg        [50:0]   ways_0_metas_22_tag;
  reg                 ways_0_metas_22_mru;
  reg                 ways_0_metas_23_vld;
  reg        [50:0]   ways_0_metas_23_tag;
  reg                 ways_0_metas_23_mru;
  reg                 ways_0_metas_24_vld;
  reg        [50:0]   ways_0_metas_24_tag;
  reg                 ways_0_metas_24_mru;
  reg                 ways_0_metas_25_vld;
  reg        [50:0]   ways_0_metas_25_tag;
  reg                 ways_0_metas_25_mru;
  reg                 ways_0_metas_26_vld;
  reg        [50:0]   ways_0_metas_26_tag;
  reg                 ways_0_metas_26_mru;
  reg                 ways_0_metas_27_vld;
  reg        [50:0]   ways_0_metas_27_tag;
  reg                 ways_0_metas_27_mru;
  reg                 ways_0_metas_28_vld;
  reg        [50:0]   ways_0_metas_28_tag;
  reg                 ways_0_metas_28_mru;
  reg                 ways_0_metas_29_vld;
  reg        [50:0]   ways_0_metas_29_tag;
  reg                 ways_0_metas_29_mru;
  reg                 ways_0_metas_30_vld;
  reg        [50:0]   ways_0_metas_30_tag;
  reg                 ways_0_metas_30_mru;
  reg                 ways_0_metas_31_vld;
  reg        [50:0]   ways_0_metas_31_tag;
  reg                 ways_0_metas_31_mru;
  reg                 ways_0_metas_32_vld;
  reg        [50:0]   ways_0_metas_32_tag;
  reg                 ways_0_metas_32_mru;
  reg                 ways_0_metas_33_vld;
  reg        [50:0]   ways_0_metas_33_tag;
  reg                 ways_0_metas_33_mru;
  reg                 ways_0_metas_34_vld;
  reg        [50:0]   ways_0_metas_34_tag;
  reg                 ways_0_metas_34_mru;
  reg                 ways_0_metas_35_vld;
  reg        [50:0]   ways_0_metas_35_tag;
  reg                 ways_0_metas_35_mru;
  reg                 ways_0_metas_36_vld;
  reg        [50:0]   ways_0_metas_36_tag;
  reg                 ways_0_metas_36_mru;
  reg                 ways_0_metas_37_vld;
  reg        [50:0]   ways_0_metas_37_tag;
  reg                 ways_0_metas_37_mru;
  reg                 ways_0_metas_38_vld;
  reg        [50:0]   ways_0_metas_38_tag;
  reg                 ways_0_metas_38_mru;
  reg                 ways_0_metas_39_vld;
  reg        [50:0]   ways_0_metas_39_tag;
  reg                 ways_0_metas_39_mru;
  reg                 ways_0_metas_40_vld;
  reg        [50:0]   ways_0_metas_40_tag;
  reg                 ways_0_metas_40_mru;
  reg                 ways_0_metas_41_vld;
  reg        [50:0]   ways_0_metas_41_tag;
  reg                 ways_0_metas_41_mru;
  reg                 ways_0_metas_42_vld;
  reg        [50:0]   ways_0_metas_42_tag;
  reg                 ways_0_metas_42_mru;
  reg                 ways_0_metas_43_vld;
  reg        [50:0]   ways_0_metas_43_tag;
  reg                 ways_0_metas_43_mru;
  reg                 ways_0_metas_44_vld;
  reg        [50:0]   ways_0_metas_44_tag;
  reg                 ways_0_metas_44_mru;
  reg                 ways_0_metas_45_vld;
  reg        [50:0]   ways_0_metas_45_tag;
  reg                 ways_0_metas_45_mru;
  reg                 ways_0_metas_46_vld;
  reg        [50:0]   ways_0_metas_46_tag;
  reg                 ways_0_metas_46_mru;
  reg                 ways_0_metas_47_vld;
  reg        [50:0]   ways_0_metas_47_tag;
  reg                 ways_0_metas_47_mru;
  reg                 ways_0_metas_48_vld;
  reg        [50:0]   ways_0_metas_48_tag;
  reg                 ways_0_metas_48_mru;
  reg                 ways_0_metas_49_vld;
  reg        [50:0]   ways_0_metas_49_tag;
  reg                 ways_0_metas_49_mru;
  reg                 ways_0_metas_50_vld;
  reg        [50:0]   ways_0_metas_50_tag;
  reg                 ways_0_metas_50_mru;
  reg                 ways_0_metas_51_vld;
  reg        [50:0]   ways_0_metas_51_tag;
  reg                 ways_0_metas_51_mru;
  reg                 ways_0_metas_52_vld;
  reg        [50:0]   ways_0_metas_52_tag;
  reg                 ways_0_metas_52_mru;
  reg                 ways_0_metas_53_vld;
  reg        [50:0]   ways_0_metas_53_tag;
  reg                 ways_0_metas_53_mru;
  reg                 ways_0_metas_54_vld;
  reg        [50:0]   ways_0_metas_54_tag;
  reg                 ways_0_metas_54_mru;
  reg                 ways_0_metas_55_vld;
  reg        [50:0]   ways_0_metas_55_tag;
  reg                 ways_0_metas_55_mru;
  reg                 ways_0_metas_56_vld;
  reg        [50:0]   ways_0_metas_56_tag;
  reg                 ways_0_metas_56_mru;
  reg                 ways_0_metas_57_vld;
  reg        [50:0]   ways_0_metas_57_tag;
  reg                 ways_0_metas_57_mru;
  reg                 ways_0_metas_58_vld;
  reg        [50:0]   ways_0_metas_58_tag;
  reg                 ways_0_metas_58_mru;
  reg                 ways_0_metas_59_vld;
  reg        [50:0]   ways_0_metas_59_tag;
  reg                 ways_0_metas_59_mru;
  reg                 ways_0_metas_60_vld;
  reg        [50:0]   ways_0_metas_60_tag;
  reg                 ways_0_metas_60_mru;
  reg                 ways_0_metas_61_vld;
  reg        [50:0]   ways_0_metas_61_tag;
  reg                 ways_0_metas_61_mru;
  reg                 ways_0_metas_62_vld;
  reg        [50:0]   ways_0_metas_62_tag;
  reg                 ways_0_metas_62_mru;
  reg                 ways_0_metas_63_vld;
  reg        [50:0]   ways_0_metas_63_tag;
  reg                 ways_0_metas_63_mru;
  reg                 ways_0_metas_64_vld;
  reg        [50:0]   ways_0_metas_64_tag;
  reg                 ways_0_metas_64_mru;
  reg                 ways_0_metas_65_vld;
  reg        [50:0]   ways_0_metas_65_tag;
  reg                 ways_0_metas_65_mru;
  reg                 ways_0_metas_66_vld;
  reg        [50:0]   ways_0_metas_66_tag;
  reg                 ways_0_metas_66_mru;
  reg                 ways_0_metas_67_vld;
  reg        [50:0]   ways_0_metas_67_tag;
  reg                 ways_0_metas_67_mru;
  reg                 ways_0_metas_68_vld;
  reg        [50:0]   ways_0_metas_68_tag;
  reg                 ways_0_metas_68_mru;
  reg                 ways_0_metas_69_vld;
  reg        [50:0]   ways_0_metas_69_tag;
  reg                 ways_0_metas_69_mru;
  reg                 ways_0_metas_70_vld;
  reg        [50:0]   ways_0_metas_70_tag;
  reg                 ways_0_metas_70_mru;
  reg                 ways_0_metas_71_vld;
  reg        [50:0]   ways_0_metas_71_tag;
  reg                 ways_0_metas_71_mru;
  reg                 ways_0_metas_72_vld;
  reg        [50:0]   ways_0_metas_72_tag;
  reg                 ways_0_metas_72_mru;
  reg                 ways_0_metas_73_vld;
  reg        [50:0]   ways_0_metas_73_tag;
  reg                 ways_0_metas_73_mru;
  reg                 ways_0_metas_74_vld;
  reg        [50:0]   ways_0_metas_74_tag;
  reg                 ways_0_metas_74_mru;
  reg                 ways_0_metas_75_vld;
  reg        [50:0]   ways_0_metas_75_tag;
  reg                 ways_0_metas_75_mru;
  reg                 ways_0_metas_76_vld;
  reg        [50:0]   ways_0_metas_76_tag;
  reg                 ways_0_metas_76_mru;
  reg                 ways_0_metas_77_vld;
  reg        [50:0]   ways_0_metas_77_tag;
  reg                 ways_0_metas_77_mru;
  reg                 ways_0_metas_78_vld;
  reg        [50:0]   ways_0_metas_78_tag;
  reg                 ways_0_metas_78_mru;
  reg                 ways_0_metas_79_vld;
  reg        [50:0]   ways_0_metas_79_tag;
  reg                 ways_0_metas_79_mru;
  reg                 ways_0_metas_80_vld;
  reg        [50:0]   ways_0_metas_80_tag;
  reg                 ways_0_metas_80_mru;
  reg                 ways_0_metas_81_vld;
  reg        [50:0]   ways_0_metas_81_tag;
  reg                 ways_0_metas_81_mru;
  reg                 ways_0_metas_82_vld;
  reg        [50:0]   ways_0_metas_82_tag;
  reg                 ways_0_metas_82_mru;
  reg                 ways_0_metas_83_vld;
  reg        [50:0]   ways_0_metas_83_tag;
  reg                 ways_0_metas_83_mru;
  reg                 ways_0_metas_84_vld;
  reg        [50:0]   ways_0_metas_84_tag;
  reg                 ways_0_metas_84_mru;
  reg                 ways_0_metas_85_vld;
  reg        [50:0]   ways_0_metas_85_tag;
  reg                 ways_0_metas_85_mru;
  reg                 ways_0_metas_86_vld;
  reg        [50:0]   ways_0_metas_86_tag;
  reg                 ways_0_metas_86_mru;
  reg                 ways_0_metas_87_vld;
  reg        [50:0]   ways_0_metas_87_tag;
  reg                 ways_0_metas_87_mru;
  reg                 ways_0_metas_88_vld;
  reg        [50:0]   ways_0_metas_88_tag;
  reg                 ways_0_metas_88_mru;
  reg                 ways_0_metas_89_vld;
  reg        [50:0]   ways_0_metas_89_tag;
  reg                 ways_0_metas_89_mru;
  reg                 ways_0_metas_90_vld;
  reg        [50:0]   ways_0_metas_90_tag;
  reg                 ways_0_metas_90_mru;
  reg                 ways_0_metas_91_vld;
  reg        [50:0]   ways_0_metas_91_tag;
  reg                 ways_0_metas_91_mru;
  reg                 ways_0_metas_92_vld;
  reg        [50:0]   ways_0_metas_92_tag;
  reg                 ways_0_metas_92_mru;
  reg                 ways_0_metas_93_vld;
  reg        [50:0]   ways_0_metas_93_tag;
  reg                 ways_0_metas_93_mru;
  reg                 ways_0_metas_94_vld;
  reg        [50:0]   ways_0_metas_94_tag;
  reg                 ways_0_metas_94_mru;
  reg                 ways_0_metas_95_vld;
  reg        [50:0]   ways_0_metas_95_tag;
  reg                 ways_0_metas_95_mru;
  reg                 ways_0_metas_96_vld;
  reg        [50:0]   ways_0_metas_96_tag;
  reg                 ways_0_metas_96_mru;
  reg                 ways_0_metas_97_vld;
  reg        [50:0]   ways_0_metas_97_tag;
  reg                 ways_0_metas_97_mru;
  reg                 ways_0_metas_98_vld;
  reg        [50:0]   ways_0_metas_98_tag;
  reg                 ways_0_metas_98_mru;
  reg                 ways_0_metas_99_vld;
  reg        [50:0]   ways_0_metas_99_tag;
  reg                 ways_0_metas_99_mru;
  reg                 ways_0_metas_100_vld;
  reg        [50:0]   ways_0_metas_100_tag;
  reg                 ways_0_metas_100_mru;
  reg                 ways_0_metas_101_vld;
  reg        [50:0]   ways_0_metas_101_tag;
  reg                 ways_0_metas_101_mru;
  reg                 ways_0_metas_102_vld;
  reg        [50:0]   ways_0_metas_102_tag;
  reg                 ways_0_metas_102_mru;
  reg                 ways_0_metas_103_vld;
  reg        [50:0]   ways_0_metas_103_tag;
  reg                 ways_0_metas_103_mru;
  reg                 ways_0_metas_104_vld;
  reg        [50:0]   ways_0_metas_104_tag;
  reg                 ways_0_metas_104_mru;
  reg                 ways_0_metas_105_vld;
  reg        [50:0]   ways_0_metas_105_tag;
  reg                 ways_0_metas_105_mru;
  reg                 ways_0_metas_106_vld;
  reg        [50:0]   ways_0_metas_106_tag;
  reg                 ways_0_metas_106_mru;
  reg                 ways_0_metas_107_vld;
  reg        [50:0]   ways_0_metas_107_tag;
  reg                 ways_0_metas_107_mru;
  reg                 ways_0_metas_108_vld;
  reg        [50:0]   ways_0_metas_108_tag;
  reg                 ways_0_metas_108_mru;
  reg                 ways_0_metas_109_vld;
  reg        [50:0]   ways_0_metas_109_tag;
  reg                 ways_0_metas_109_mru;
  reg                 ways_0_metas_110_vld;
  reg        [50:0]   ways_0_metas_110_tag;
  reg                 ways_0_metas_110_mru;
  reg                 ways_0_metas_111_vld;
  reg        [50:0]   ways_0_metas_111_tag;
  reg                 ways_0_metas_111_mru;
  reg                 ways_0_metas_112_vld;
  reg        [50:0]   ways_0_metas_112_tag;
  reg                 ways_0_metas_112_mru;
  reg                 ways_0_metas_113_vld;
  reg        [50:0]   ways_0_metas_113_tag;
  reg                 ways_0_metas_113_mru;
  reg                 ways_0_metas_114_vld;
  reg        [50:0]   ways_0_metas_114_tag;
  reg                 ways_0_metas_114_mru;
  reg                 ways_0_metas_115_vld;
  reg        [50:0]   ways_0_metas_115_tag;
  reg                 ways_0_metas_115_mru;
  reg                 ways_0_metas_116_vld;
  reg        [50:0]   ways_0_metas_116_tag;
  reg                 ways_0_metas_116_mru;
  reg                 ways_0_metas_117_vld;
  reg        [50:0]   ways_0_metas_117_tag;
  reg                 ways_0_metas_117_mru;
  reg                 ways_0_metas_118_vld;
  reg        [50:0]   ways_0_metas_118_tag;
  reg                 ways_0_metas_118_mru;
  reg                 ways_0_metas_119_vld;
  reg        [50:0]   ways_0_metas_119_tag;
  reg                 ways_0_metas_119_mru;
  reg                 ways_0_metas_120_vld;
  reg        [50:0]   ways_0_metas_120_tag;
  reg                 ways_0_metas_120_mru;
  reg                 ways_0_metas_121_vld;
  reg        [50:0]   ways_0_metas_121_tag;
  reg                 ways_0_metas_121_mru;
  reg                 ways_0_metas_122_vld;
  reg        [50:0]   ways_0_metas_122_tag;
  reg                 ways_0_metas_122_mru;
  reg                 ways_0_metas_123_vld;
  reg        [50:0]   ways_0_metas_123_tag;
  reg                 ways_0_metas_123_mru;
  reg                 ways_0_metas_124_vld;
  reg        [50:0]   ways_0_metas_124_tag;
  reg                 ways_0_metas_124_mru;
  reg                 ways_0_metas_125_vld;
  reg        [50:0]   ways_0_metas_125_tag;
  reg                 ways_0_metas_125_mru;
  reg                 ways_0_metas_126_vld;
  reg        [50:0]   ways_0_metas_126_tag;
  reg                 ways_0_metas_126_mru;
  reg                 ways_0_metas_127_vld;
  reg        [50:0]   ways_0_metas_127_tag;
  reg                 ways_0_metas_127_mru;
  reg                 ways_1_metas_0_vld;
  reg        [50:0]   ways_1_metas_0_tag;
  reg                 ways_1_metas_0_mru;
  reg                 ways_1_metas_1_vld;
  reg        [50:0]   ways_1_metas_1_tag;
  reg                 ways_1_metas_1_mru;
  reg                 ways_1_metas_2_vld;
  reg        [50:0]   ways_1_metas_2_tag;
  reg                 ways_1_metas_2_mru;
  reg                 ways_1_metas_3_vld;
  reg        [50:0]   ways_1_metas_3_tag;
  reg                 ways_1_metas_3_mru;
  reg                 ways_1_metas_4_vld;
  reg        [50:0]   ways_1_metas_4_tag;
  reg                 ways_1_metas_4_mru;
  reg                 ways_1_metas_5_vld;
  reg        [50:0]   ways_1_metas_5_tag;
  reg                 ways_1_metas_5_mru;
  reg                 ways_1_metas_6_vld;
  reg        [50:0]   ways_1_metas_6_tag;
  reg                 ways_1_metas_6_mru;
  reg                 ways_1_metas_7_vld;
  reg        [50:0]   ways_1_metas_7_tag;
  reg                 ways_1_metas_7_mru;
  reg                 ways_1_metas_8_vld;
  reg        [50:0]   ways_1_metas_8_tag;
  reg                 ways_1_metas_8_mru;
  reg                 ways_1_metas_9_vld;
  reg        [50:0]   ways_1_metas_9_tag;
  reg                 ways_1_metas_9_mru;
  reg                 ways_1_metas_10_vld;
  reg        [50:0]   ways_1_metas_10_tag;
  reg                 ways_1_metas_10_mru;
  reg                 ways_1_metas_11_vld;
  reg        [50:0]   ways_1_metas_11_tag;
  reg                 ways_1_metas_11_mru;
  reg                 ways_1_metas_12_vld;
  reg        [50:0]   ways_1_metas_12_tag;
  reg                 ways_1_metas_12_mru;
  reg                 ways_1_metas_13_vld;
  reg        [50:0]   ways_1_metas_13_tag;
  reg                 ways_1_metas_13_mru;
  reg                 ways_1_metas_14_vld;
  reg        [50:0]   ways_1_metas_14_tag;
  reg                 ways_1_metas_14_mru;
  reg                 ways_1_metas_15_vld;
  reg        [50:0]   ways_1_metas_15_tag;
  reg                 ways_1_metas_15_mru;
  reg                 ways_1_metas_16_vld;
  reg        [50:0]   ways_1_metas_16_tag;
  reg                 ways_1_metas_16_mru;
  reg                 ways_1_metas_17_vld;
  reg        [50:0]   ways_1_metas_17_tag;
  reg                 ways_1_metas_17_mru;
  reg                 ways_1_metas_18_vld;
  reg        [50:0]   ways_1_metas_18_tag;
  reg                 ways_1_metas_18_mru;
  reg                 ways_1_metas_19_vld;
  reg        [50:0]   ways_1_metas_19_tag;
  reg                 ways_1_metas_19_mru;
  reg                 ways_1_metas_20_vld;
  reg        [50:0]   ways_1_metas_20_tag;
  reg                 ways_1_metas_20_mru;
  reg                 ways_1_metas_21_vld;
  reg        [50:0]   ways_1_metas_21_tag;
  reg                 ways_1_metas_21_mru;
  reg                 ways_1_metas_22_vld;
  reg        [50:0]   ways_1_metas_22_tag;
  reg                 ways_1_metas_22_mru;
  reg                 ways_1_metas_23_vld;
  reg        [50:0]   ways_1_metas_23_tag;
  reg                 ways_1_metas_23_mru;
  reg                 ways_1_metas_24_vld;
  reg        [50:0]   ways_1_metas_24_tag;
  reg                 ways_1_metas_24_mru;
  reg                 ways_1_metas_25_vld;
  reg        [50:0]   ways_1_metas_25_tag;
  reg                 ways_1_metas_25_mru;
  reg                 ways_1_metas_26_vld;
  reg        [50:0]   ways_1_metas_26_tag;
  reg                 ways_1_metas_26_mru;
  reg                 ways_1_metas_27_vld;
  reg        [50:0]   ways_1_metas_27_tag;
  reg                 ways_1_metas_27_mru;
  reg                 ways_1_metas_28_vld;
  reg        [50:0]   ways_1_metas_28_tag;
  reg                 ways_1_metas_28_mru;
  reg                 ways_1_metas_29_vld;
  reg        [50:0]   ways_1_metas_29_tag;
  reg                 ways_1_metas_29_mru;
  reg                 ways_1_metas_30_vld;
  reg        [50:0]   ways_1_metas_30_tag;
  reg                 ways_1_metas_30_mru;
  reg                 ways_1_metas_31_vld;
  reg        [50:0]   ways_1_metas_31_tag;
  reg                 ways_1_metas_31_mru;
  reg                 ways_1_metas_32_vld;
  reg        [50:0]   ways_1_metas_32_tag;
  reg                 ways_1_metas_32_mru;
  reg                 ways_1_metas_33_vld;
  reg        [50:0]   ways_1_metas_33_tag;
  reg                 ways_1_metas_33_mru;
  reg                 ways_1_metas_34_vld;
  reg        [50:0]   ways_1_metas_34_tag;
  reg                 ways_1_metas_34_mru;
  reg                 ways_1_metas_35_vld;
  reg        [50:0]   ways_1_metas_35_tag;
  reg                 ways_1_metas_35_mru;
  reg                 ways_1_metas_36_vld;
  reg        [50:0]   ways_1_metas_36_tag;
  reg                 ways_1_metas_36_mru;
  reg                 ways_1_metas_37_vld;
  reg        [50:0]   ways_1_metas_37_tag;
  reg                 ways_1_metas_37_mru;
  reg                 ways_1_metas_38_vld;
  reg        [50:0]   ways_1_metas_38_tag;
  reg                 ways_1_metas_38_mru;
  reg                 ways_1_metas_39_vld;
  reg        [50:0]   ways_1_metas_39_tag;
  reg                 ways_1_metas_39_mru;
  reg                 ways_1_metas_40_vld;
  reg        [50:0]   ways_1_metas_40_tag;
  reg                 ways_1_metas_40_mru;
  reg                 ways_1_metas_41_vld;
  reg        [50:0]   ways_1_metas_41_tag;
  reg                 ways_1_metas_41_mru;
  reg                 ways_1_metas_42_vld;
  reg        [50:0]   ways_1_metas_42_tag;
  reg                 ways_1_metas_42_mru;
  reg                 ways_1_metas_43_vld;
  reg        [50:0]   ways_1_metas_43_tag;
  reg                 ways_1_metas_43_mru;
  reg                 ways_1_metas_44_vld;
  reg        [50:0]   ways_1_metas_44_tag;
  reg                 ways_1_metas_44_mru;
  reg                 ways_1_metas_45_vld;
  reg        [50:0]   ways_1_metas_45_tag;
  reg                 ways_1_metas_45_mru;
  reg                 ways_1_metas_46_vld;
  reg        [50:0]   ways_1_metas_46_tag;
  reg                 ways_1_metas_46_mru;
  reg                 ways_1_metas_47_vld;
  reg        [50:0]   ways_1_metas_47_tag;
  reg                 ways_1_metas_47_mru;
  reg                 ways_1_metas_48_vld;
  reg        [50:0]   ways_1_metas_48_tag;
  reg                 ways_1_metas_48_mru;
  reg                 ways_1_metas_49_vld;
  reg        [50:0]   ways_1_metas_49_tag;
  reg                 ways_1_metas_49_mru;
  reg                 ways_1_metas_50_vld;
  reg        [50:0]   ways_1_metas_50_tag;
  reg                 ways_1_metas_50_mru;
  reg                 ways_1_metas_51_vld;
  reg        [50:0]   ways_1_metas_51_tag;
  reg                 ways_1_metas_51_mru;
  reg                 ways_1_metas_52_vld;
  reg        [50:0]   ways_1_metas_52_tag;
  reg                 ways_1_metas_52_mru;
  reg                 ways_1_metas_53_vld;
  reg        [50:0]   ways_1_metas_53_tag;
  reg                 ways_1_metas_53_mru;
  reg                 ways_1_metas_54_vld;
  reg        [50:0]   ways_1_metas_54_tag;
  reg                 ways_1_metas_54_mru;
  reg                 ways_1_metas_55_vld;
  reg        [50:0]   ways_1_metas_55_tag;
  reg                 ways_1_metas_55_mru;
  reg                 ways_1_metas_56_vld;
  reg        [50:0]   ways_1_metas_56_tag;
  reg                 ways_1_metas_56_mru;
  reg                 ways_1_metas_57_vld;
  reg        [50:0]   ways_1_metas_57_tag;
  reg                 ways_1_metas_57_mru;
  reg                 ways_1_metas_58_vld;
  reg        [50:0]   ways_1_metas_58_tag;
  reg                 ways_1_metas_58_mru;
  reg                 ways_1_metas_59_vld;
  reg        [50:0]   ways_1_metas_59_tag;
  reg                 ways_1_metas_59_mru;
  reg                 ways_1_metas_60_vld;
  reg        [50:0]   ways_1_metas_60_tag;
  reg                 ways_1_metas_60_mru;
  reg                 ways_1_metas_61_vld;
  reg        [50:0]   ways_1_metas_61_tag;
  reg                 ways_1_metas_61_mru;
  reg                 ways_1_metas_62_vld;
  reg        [50:0]   ways_1_metas_62_tag;
  reg                 ways_1_metas_62_mru;
  reg                 ways_1_metas_63_vld;
  reg        [50:0]   ways_1_metas_63_tag;
  reg                 ways_1_metas_63_mru;
  reg                 ways_1_metas_64_vld;
  reg        [50:0]   ways_1_metas_64_tag;
  reg                 ways_1_metas_64_mru;
  reg                 ways_1_metas_65_vld;
  reg        [50:0]   ways_1_metas_65_tag;
  reg                 ways_1_metas_65_mru;
  reg                 ways_1_metas_66_vld;
  reg        [50:0]   ways_1_metas_66_tag;
  reg                 ways_1_metas_66_mru;
  reg                 ways_1_metas_67_vld;
  reg        [50:0]   ways_1_metas_67_tag;
  reg                 ways_1_metas_67_mru;
  reg                 ways_1_metas_68_vld;
  reg        [50:0]   ways_1_metas_68_tag;
  reg                 ways_1_metas_68_mru;
  reg                 ways_1_metas_69_vld;
  reg        [50:0]   ways_1_metas_69_tag;
  reg                 ways_1_metas_69_mru;
  reg                 ways_1_metas_70_vld;
  reg        [50:0]   ways_1_metas_70_tag;
  reg                 ways_1_metas_70_mru;
  reg                 ways_1_metas_71_vld;
  reg        [50:0]   ways_1_metas_71_tag;
  reg                 ways_1_metas_71_mru;
  reg                 ways_1_metas_72_vld;
  reg        [50:0]   ways_1_metas_72_tag;
  reg                 ways_1_metas_72_mru;
  reg                 ways_1_metas_73_vld;
  reg        [50:0]   ways_1_metas_73_tag;
  reg                 ways_1_metas_73_mru;
  reg                 ways_1_metas_74_vld;
  reg        [50:0]   ways_1_metas_74_tag;
  reg                 ways_1_metas_74_mru;
  reg                 ways_1_metas_75_vld;
  reg        [50:0]   ways_1_metas_75_tag;
  reg                 ways_1_metas_75_mru;
  reg                 ways_1_metas_76_vld;
  reg        [50:0]   ways_1_metas_76_tag;
  reg                 ways_1_metas_76_mru;
  reg                 ways_1_metas_77_vld;
  reg        [50:0]   ways_1_metas_77_tag;
  reg                 ways_1_metas_77_mru;
  reg                 ways_1_metas_78_vld;
  reg        [50:0]   ways_1_metas_78_tag;
  reg                 ways_1_metas_78_mru;
  reg                 ways_1_metas_79_vld;
  reg        [50:0]   ways_1_metas_79_tag;
  reg                 ways_1_metas_79_mru;
  reg                 ways_1_metas_80_vld;
  reg        [50:0]   ways_1_metas_80_tag;
  reg                 ways_1_metas_80_mru;
  reg                 ways_1_metas_81_vld;
  reg        [50:0]   ways_1_metas_81_tag;
  reg                 ways_1_metas_81_mru;
  reg                 ways_1_metas_82_vld;
  reg        [50:0]   ways_1_metas_82_tag;
  reg                 ways_1_metas_82_mru;
  reg                 ways_1_metas_83_vld;
  reg        [50:0]   ways_1_metas_83_tag;
  reg                 ways_1_metas_83_mru;
  reg                 ways_1_metas_84_vld;
  reg        [50:0]   ways_1_metas_84_tag;
  reg                 ways_1_metas_84_mru;
  reg                 ways_1_metas_85_vld;
  reg        [50:0]   ways_1_metas_85_tag;
  reg                 ways_1_metas_85_mru;
  reg                 ways_1_metas_86_vld;
  reg        [50:0]   ways_1_metas_86_tag;
  reg                 ways_1_metas_86_mru;
  reg                 ways_1_metas_87_vld;
  reg        [50:0]   ways_1_metas_87_tag;
  reg                 ways_1_metas_87_mru;
  reg                 ways_1_metas_88_vld;
  reg        [50:0]   ways_1_metas_88_tag;
  reg                 ways_1_metas_88_mru;
  reg                 ways_1_metas_89_vld;
  reg        [50:0]   ways_1_metas_89_tag;
  reg                 ways_1_metas_89_mru;
  reg                 ways_1_metas_90_vld;
  reg        [50:0]   ways_1_metas_90_tag;
  reg                 ways_1_metas_90_mru;
  reg                 ways_1_metas_91_vld;
  reg        [50:0]   ways_1_metas_91_tag;
  reg                 ways_1_metas_91_mru;
  reg                 ways_1_metas_92_vld;
  reg        [50:0]   ways_1_metas_92_tag;
  reg                 ways_1_metas_92_mru;
  reg                 ways_1_metas_93_vld;
  reg        [50:0]   ways_1_metas_93_tag;
  reg                 ways_1_metas_93_mru;
  reg                 ways_1_metas_94_vld;
  reg        [50:0]   ways_1_metas_94_tag;
  reg                 ways_1_metas_94_mru;
  reg                 ways_1_metas_95_vld;
  reg        [50:0]   ways_1_metas_95_tag;
  reg                 ways_1_metas_95_mru;
  reg                 ways_1_metas_96_vld;
  reg        [50:0]   ways_1_metas_96_tag;
  reg                 ways_1_metas_96_mru;
  reg                 ways_1_metas_97_vld;
  reg        [50:0]   ways_1_metas_97_tag;
  reg                 ways_1_metas_97_mru;
  reg                 ways_1_metas_98_vld;
  reg        [50:0]   ways_1_metas_98_tag;
  reg                 ways_1_metas_98_mru;
  reg                 ways_1_metas_99_vld;
  reg        [50:0]   ways_1_metas_99_tag;
  reg                 ways_1_metas_99_mru;
  reg                 ways_1_metas_100_vld;
  reg        [50:0]   ways_1_metas_100_tag;
  reg                 ways_1_metas_100_mru;
  reg                 ways_1_metas_101_vld;
  reg        [50:0]   ways_1_metas_101_tag;
  reg                 ways_1_metas_101_mru;
  reg                 ways_1_metas_102_vld;
  reg        [50:0]   ways_1_metas_102_tag;
  reg                 ways_1_metas_102_mru;
  reg                 ways_1_metas_103_vld;
  reg        [50:0]   ways_1_metas_103_tag;
  reg                 ways_1_metas_103_mru;
  reg                 ways_1_metas_104_vld;
  reg        [50:0]   ways_1_metas_104_tag;
  reg                 ways_1_metas_104_mru;
  reg                 ways_1_metas_105_vld;
  reg        [50:0]   ways_1_metas_105_tag;
  reg                 ways_1_metas_105_mru;
  reg                 ways_1_metas_106_vld;
  reg        [50:0]   ways_1_metas_106_tag;
  reg                 ways_1_metas_106_mru;
  reg                 ways_1_metas_107_vld;
  reg        [50:0]   ways_1_metas_107_tag;
  reg                 ways_1_metas_107_mru;
  reg                 ways_1_metas_108_vld;
  reg        [50:0]   ways_1_metas_108_tag;
  reg                 ways_1_metas_108_mru;
  reg                 ways_1_metas_109_vld;
  reg        [50:0]   ways_1_metas_109_tag;
  reg                 ways_1_metas_109_mru;
  reg                 ways_1_metas_110_vld;
  reg        [50:0]   ways_1_metas_110_tag;
  reg                 ways_1_metas_110_mru;
  reg                 ways_1_metas_111_vld;
  reg        [50:0]   ways_1_metas_111_tag;
  reg                 ways_1_metas_111_mru;
  reg                 ways_1_metas_112_vld;
  reg        [50:0]   ways_1_metas_112_tag;
  reg                 ways_1_metas_112_mru;
  reg                 ways_1_metas_113_vld;
  reg        [50:0]   ways_1_metas_113_tag;
  reg                 ways_1_metas_113_mru;
  reg                 ways_1_metas_114_vld;
  reg        [50:0]   ways_1_metas_114_tag;
  reg                 ways_1_metas_114_mru;
  reg                 ways_1_metas_115_vld;
  reg        [50:0]   ways_1_metas_115_tag;
  reg                 ways_1_metas_115_mru;
  reg                 ways_1_metas_116_vld;
  reg        [50:0]   ways_1_metas_116_tag;
  reg                 ways_1_metas_116_mru;
  reg                 ways_1_metas_117_vld;
  reg        [50:0]   ways_1_metas_117_tag;
  reg                 ways_1_metas_117_mru;
  reg                 ways_1_metas_118_vld;
  reg        [50:0]   ways_1_metas_118_tag;
  reg                 ways_1_metas_118_mru;
  reg                 ways_1_metas_119_vld;
  reg        [50:0]   ways_1_metas_119_tag;
  reg                 ways_1_metas_119_mru;
  reg                 ways_1_metas_120_vld;
  reg        [50:0]   ways_1_metas_120_tag;
  reg                 ways_1_metas_120_mru;
  reg                 ways_1_metas_121_vld;
  reg        [50:0]   ways_1_metas_121_tag;
  reg                 ways_1_metas_121_mru;
  reg                 ways_1_metas_122_vld;
  reg        [50:0]   ways_1_metas_122_tag;
  reg                 ways_1_metas_122_mru;
  reg                 ways_1_metas_123_vld;
  reg        [50:0]   ways_1_metas_123_tag;
  reg                 ways_1_metas_123_mru;
  reg                 ways_1_metas_124_vld;
  reg        [50:0]   ways_1_metas_124_tag;
  reg                 ways_1_metas_124_mru;
  reg                 ways_1_metas_125_vld;
  reg        [50:0]   ways_1_metas_125_tag;
  reg                 ways_1_metas_125_mru;
  reg                 ways_1_metas_126_vld;
  reg        [50:0]   ways_1_metas_126_tag;
  reg                 ways_1_metas_126_mru;
  reg                 ways_1_metas_127_vld;
  reg        [50:0]   ways_1_metas_127_tag;
  reg                 ways_1_metas_127_mru;
  reg                 ways_2_metas_0_vld;
  reg        [50:0]   ways_2_metas_0_tag;
  reg                 ways_2_metas_0_mru;
  reg                 ways_2_metas_1_vld;
  reg        [50:0]   ways_2_metas_1_tag;
  reg                 ways_2_metas_1_mru;
  reg                 ways_2_metas_2_vld;
  reg        [50:0]   ways_2_metas_2_tag;
  reg                 ways_2_metas_2_mru;
  reg                 ways_2_metas_3_vld;
  reg        [50:0]   ways_2_metas_3_tag;
  reg                 ways_2_metas_3_mru;
  reg                 ways_2_metas_4_vld;
  reg        [50:0]   ways_2_metas_4_tag;
  reg                 ways_2_metas_4_mru;
  reg                 ways_2_metas_5_vld;
  reg        [50:0]   ways_2_metas_5_tag;
  reg                 ways_2_metas_5_mru;
  reg                 ways_2_metas_6_vld;
  reg        [50:0]   ways_2_metas_6_tag;
  reg                 ways_2_metas_6_mru;
  reg                 ways_2_metas_7_vld;
  reg        [50:0]   ways_2_metas_7_tag;
  reg                 ways_2_metas_7_mru;
  reg                 ways_2_metas_8_vld;
  reg        [50:0]   ways_2_metas_8_tag;
  reg                 ways_2_metas_8_mru;
  reg                 ways_2_metas_9_vld;
  reg        [50:0]   ways_2_metas_9_tag;
  reg                 ways_2_metas_9_mru;
  reg                 ways_2_metas_10_vld;
  reg        [50:0]   ways_2_metas_10_tag;
  reg                 ways_2_metas_10_mru;
  reg                 ways_2_metas_11_vld;
  reg        [50:0]   ways_2_metas_11_tag;
  reg                 ways_2_metas_11_mru;
  reg                 ways_2_metas_12_vld;
  reg        [50:0]   ways_2_metas_12_tag;
  reg                 ways_2_metas_12_mru;
  reg                 ways_2_metas_13_vld;
  reg        [50:0]   ways_2_metas_13_tag;
  reg                 ways_2_metas_13_mru;
  reg                 ways_2_metas_14_vld;
  reg        [50:0]   ways_2_metas_14_tag;
  reg                 ways_2_metas_14_mru;
  reg                 ways_2_metas_15_vld;
  reg        [50:0]   ways_2_metas_15_tag;
  reg                 ways_2_metas_15_mru;
  reg                 ways_2_metas_16_vld;
  reg        [50:0]   ways_2_metas_16_tag;
  reg                 ways_2_metas_16_mru;
  reg                 ways_2_metas_17_vld;
  reg        [50:0]   ways_2_metas_17_tag;
  reg                 ways_2_metas_17_mru;
  reg                 ways_2_metas_18_vld;
  reg        [50:0]   ways_2_metas_18_tag;
  reg                 ways_2_metas_18_mru;
  reg                 ways_2_metas_19_vld;
  reg        [50:0]   ways_2_metas_19_tag;
  reg                 ways_2_metas_19_mru;
  reg                 ways_2_metas_20_vld;
  reg        [50:0]   ways_2_metas_20_tag;
  reg                 ways_2_metas_20_mru;
  reg                 ways_2_metas_21_vld;
  reg        [50:0]   ways_2_metas_21_tag;
  reg                 ways_2_metas_21_mru;
  reg                 ways_2_metas_22_vld;
  reg        [50:0]   ways_2_metas_22_tag;
  reg                 ways_2_metas_22_mru;
  reg                 ways_2_metas_23_vld;
  reg        [50:0]   ways_2_metas_23_tag;
  reg                 ways_2_metas_23_mru;
  reg                 ways_2_metas_24_vld;
  reg        [50:0]   ways_2_metas_24_tag;
  reg                 ways_2_metas_24_mru;
  reg                 ways_2_metas_25_vld;
  reg        [50:0]   ways_2_metas_25_tag;
  reg                 ways_2_metas_25_mru;
  reg                 ways_2_metas_26_vld;
  reg        [50:0]   ways_2_metas_26_tag;
  reg                 ways_2_metas_26_mru;
  reg                 ways_2_metas_27_vld;
  reg        [50:0]   ways_2_metas_27_tag;
  reg                 ways_2_metas_27_mru;
  reg                 ways_2_metas_28_vld;
  reg        [50:0]   ways_2_metas_28_tag;
  reg                 ways_2_metas_28_mru;
  reg                 ways_2_metas_29_vld;
  reg        [50:0]   ways_2_metas_29_tag;
  reg                 ways_2_metas_29_mru;
  reg                 ways_2_metas_30_vld;
  reg        [50:0]   ways_2_metas_30_tag;
  reg                 ways_2_metas_30_mru;
  reg                 ways_2_metas_31_vld;
  reg        [50:0]   ways_2_metas_31_tag;
  reg                 ways_2_metas_31_mru;
  reg                 ways_2_metas_32_vld;
  reg        [50:0]   ways_2_metas_32_tag;
  reg                 ways_2_metas_32_mru;
  reg                 ways_2_metas_33_vld;
  reg        [50:0]   ways_2_metas_33_tag;
  reg                 ways_2_metas_33_mru;
  reg                 ways_2_metas_34_vld;
  reg        [50:0]   ways_2_metas_34_tag;
  reg                 ways_2_metas_34_mru;
  reg                 ways_2_metas_35_vld;
  reg        [50:0]   ways_2_metas_35_tag;
  reg                 ways_2_metas_35_mru;
  reg                 ways_2_metas_36_vld;
  reg        [50:0]   ways_2_metas_36_tag;
  reg                 ways_2_metas_36_mru;
  reg                 ways_2_metas_37_vld;
  reg        [50:0]   ways_2_metas_37_tag;
  reg                 ways_2_metas_37_mru;
  reg                 ways_2_metas_38_vld;
  reg        [50:0]   ways_2_metas_38_tag;
  reg                 ways_2_metas_38_mru;
  reg                 ways_2_metas_39_vld;
  reg        [50:0]   ways_2_metas_39_tag;
  reg                 ways_2_metas_39_mru;
  reg                 ways_2_metas_40_vld;
  reg        [50:0]   ways_2_metas_40_tag;
  reg                 ways_2_metas_40_mru;
  reg                 ways_2_metas_41_vld;
  reg        [50:0]   ways_2_metas_41_tag;
  reg                 ways_2_metas_41_mru;
  reg                 ways_2_metas_42_vld;
  reg        [50:0]   ways_2_metas_42_tag;
  reg                 ways_2_metas_42_mru;
  reg                 ways_2_metas_43_vld;
  reg        [50:0]   ways_2_metas_43_tag;
  reg                 ways_2_metas_43_mru;
  reg                 ways_2_metas_44_vld;
  reg        [50:0]   ways_2_metas_44_tag;
  reg                 ways_2_metas_44_mru;
  reg                 ways_2_metas_45_vld;
  reg        [50:0]   ways_2_metas_45_tag;
  reg                 ways_2_metas_45_mru;
  reg                 ways_2_metas_46_vld;
  reg        [50:0]   ways_2_metas_46_tag;
  reg                 ways_2_metas_46_mru;
  reg                 ways_2_metas_47_vld;
  reg        [50:0]   ways_2_metas_47_tag;
  reg                 ways_2_metas_47_mru;
  reg                 ways_2_metas_48_vld;
  reg        [50:0]   ways_2_metas_48_tag;
  reg                 ways_2_metas_48_mru;
  reg                 ways_2_metas_49_vld;
  reg        [50:0]   ways_2_metas_49_tag;
  reg                 ways_2_metas_49_mru;
  reg                 ways_2_metas_50_vld;
  reg        [50:0]   ways_2_metas_50_tag;
  reg                 ways_2_metas_50_mru;
  reg                 ways_2_metas_51_vld;
  reg        [50:0]   ways_2_metas_51_tag;
  reg                 ways_2_metas_51_mru;
  reg                 ways_2_metas_52_vld;
  reg        [50:0]   ways_2_metas_52_tag;
  reg                 ways_2_metas_52_mru;
  reg                 ways_2_metas_53_vld;
  reg        [50:0]   ways_2_metas_53_tag;
  reg                 ways_2_metas_53_mru;
  reg                 ways_2_metas_54_vld;
  reg        [50:0]   ways_2_metas_54_tag;
  reg                 ways_2_metas_54_mru;
  reg                 ways_2_metas_55_vld;
  reg        [50:0]   ways_2_metas_55_tag;
  reg                 ways_2_metas_55_mru;
  reg                 ways_2_metas_56_vld;
  reg        [50:0]   ways_2_metas_56_tag;
  reg                 ways_2_metas_56_mru;
  reg                 ways_2_metas_57_vld;
  reg        [50:0]   ways_2_metas_57_tag;
  reg                 ways_2_metas_57_mru;
  reg                 ways_2_metas_58_vld;
  reg        [50:0]   ways_2_metas_58_tag;
  reg                 ways_2_metas_58_mru;
  reg                 ways_2_metas_59_vld;
  reg        [50:0]   ways_2_metas_59_tag;
  reg                 ways_2_metas_59_mru;
  reg                 ways_2_metas_60_vld;
  reg        [50:0]   ways_2_metas_60_tag;
  reg                 ways_2_metas_60_mru;
  reg                 ways_2_metas_61_vld;
  reg        [50:0]   ways_2_metas_61_tag;
  reg                 ways_2_metas_61_mru;
  reg                 ways_2_metas_62_vld;
  reg        [50:0]   ways_2_metas_62_tag;
  reg                 ways_2_metas_62_mru;
  reg                 ways_2_metas_63_vld;
  reg        [50:0]   ways_2_metas_63_tag;
  reg                 ways_2_metas_63_mru;
  reg                 ways_2_metas_64_vld;
  reg        [50:0]   ways_2_metas_64_tag;
  reg                 ways_2_metas_64_mru;
  reg                 ways_2_metas_65_vld;
  reg        [50:0]   ways_2_metas_65_tag;
  reg                 ways_2_metas_65_mru;
  reg                 ways_2_metas_66_vld;
  reg        [50:0]   ways_2_metas_66_tag;
  reg                 ways_2_metas_66_mru;
  reg                 ways_2_metas_67_vld;
  reg        [50:0]   ways_2_metas_67_tag;
  reg                 ways_2_metas_67_mru;
  reg                 ways_2_metas_68_vld;
  reg        [50:0]   ways_2_metas_68_tag;
  reg                 ways_2_metas_68_mru;
  reg                 ways_2_metas_69_vld;
  reg        [50:0]   ways_2_metas_69_tag;
  reg                 ways_2_metas_69_mru;
  reg                 ways_2_metas_70_vld;
  reg        [50:0]   ways_2_metas_70_tag;
  reg                 ways_2_metas_70_mru;
  reg                 ways_2_metas_71_vld;
  reg        [50:0]   ways_2_metas_71_tag;
  reg                 ways_2_metas_71_mru;
  reg                 ways_2_metas_72_vld;
  reg        [50:0]   ways_2_metas_72_tag;
  reg                 ways_2_metas_72_mru;
  reg                 ways_2_metas_73_vld;
  reg        [50:0]   ways_2_metas_73_tag;
  reg                 ways_2_metas_73_mru;
  reg                 ways_2_metas_74_vld;
  reg        [50:0]   ways_2_metas_74_tag;
  reg                 ways_2_metas_74_mru;
  reg                 ways_2_metas_75_vld;
  reg        [50:0]   ways_2_metas_75_tag;
  reg                 ways_2_metas_75_mru;
  reg                 ways_2_metas_76_vld;
  reg        [50:0]   ways_2_metas_76_tag;
  reg                 ways_2_metas_76_mru;
  reg                 ways_2_metas_77_vld;
  reg        [50:0]   ways_2_metas_77_tag;
  reg                 ways_2_metas_77_mru;
  reg                 ways_2_metas_78_vld;
  reg        [50:0]   ways_2_metas_78_tag;
  reg                 ways_2_metas_78_mru;
  reg                 ways_2_metas_79_vld;
  reg        [50:0]   ways_2_metas_79_tag;
  reg                 ways_2_metas_79_mru;
  reg                 ways_2_metas_80_vld;
  reg        [50:0]   ways_2_metas_80_tag;
  reg                 ways_2_metas_80_mru;
  reg                 ways_2_metas_81_vld;
  reg        [50:0]   ways_2_metas_81_tag;
  reg                 ways_2_metas_81_mru;
  reg                 ways_2_metas_82_vld;
  reg        [50:0]   ways_2_metas_82_tag;
  reg                 ways_2_metas_82_mru;
  reg                 ways_2_metas_83_vld;
  reg        [50:0]   ways_2_metas_83_tag;
  reg                 ways_2_metas_83_mru;
  reg                 ways_2_metas_84_vld;
  reg        [50:0]   ways_2_metas_84_tag;
  reg                 ways_2_metas_84_mru;
  reg                 ways_2_metas_85_vld;
  reg        [50:0]   ways_2_metas_85_tag;
  reg                 ways_2_metas_85_mru;
  reg                 ways_2_metas_86_vld;
  reg        [50:0]   ways_2_metas_86_tag;
  reg                 ways_2_metas_86_mru;
  reg                 ways_2_metas_87_vld;
  reg        [50:0]   ways_2_metas_87_tag;
  reg                 ways_2_metas_87_mru;
  reg                 ways_2_metas_88_vld;
  reg        [50:0]   ways_2_metas_88_tag;
  reg                 ways_2_metas_88_mru;
  reg                 ways_2_metas_89_vld;
  reg        [50:0]   ways_2_metas_89_tag;
  reg                 ways_2_metas_89_mru;
  reg                 ways_2_metas_90_vld;
  reg        [50:0]   ways_2_metas_90_tag;
  reg                 ways_2_metas_90_mru;
  reg                 ways_2_metas_91_vld;
  reg        [50:0]   ways_2_metas_91_tag;
  reg                 ways_2_metas_91_mru;
  reg                 ways_2_metas_92_vld;
  reg        [50:0]   ways_2_metas_92_tag;
  reg                 ways_2_metas_92_mru;
  reg                 ways_2_metas_93_vld;
  reg        [50:0]   ways_2_metas_93_tag;
  reg                 ways_2_metas_93_mru;
  reg                 ways_2_metas_94_vld;
  reg        [50:0]   ways_2_metas_94_tag;
  reg                 ways_2_metas_94_mru;
  reg                 ways_2_metas_95_vld;
  reg        [50:0]   ways_2_metas_95_tag;
  reg                 ways_2_metas_95_mru;
  reg                 ways_2_metas_96_vld;
  reg        [50:0]   ways_2_metas_96_tag;
  reg                 ways_2_metas_96_mru;
  reg                 ways_2_metas_97_vld;
  reg        [50:0]   ways_2_metas_97_tag;
  reg                 ways_2_metas_97_mru;
  reg                 ways_2_metas_98_vld;
  reg        [50:0]   ways_2_metas_98_tag;
  reg                 ways_2_metas_98_mru;
  reg                 ways_2_metas_99_vld;
  reg        [50:0]   ways_2_metas_99_tag;
  reg                 ways_2_metas_99_mru;
  reg                 ways_2_metas_100_vld;
  reg        [50:0]   ways_2_metas_100_tag;
  reg                 ways_2_metas_100_mru;
  reg                 ways_2_metas_101_vld;
  reg        [50:0]   ways_2_metas_101_tag;
  reg                 ways_2_metas_101_mru;
  reg                 ways_2_metas_102_vld;
  reg        [50:0]   ways_2_metas_102_tag;
  reg                 ways_2_metas_102_mru;
  reg                 ways_2_metas_103_vld;
  reg        [50:0]   ways_2_metas_103_tag;
  reg                 ways_2_metas_103_mru;
  reg                 ways_2_metas_104_vld;
  reg        [50:0]   ways_2_metas_104_tag;
  reg                 ways_2_metas_104_mru;
  reg                 ways_2_metas_105_vld;
  reg        [50:0]   ways_2_metas_105_tag;
  reg                 ways_2_metas_105_mru;
  reg                 ways_2_metas_106_vld;
  reg        [50:0]   ways_2_metas_106_tag;
  reg                 ways_2_metas_106_mru;
  reg                 ways_2_metas_107_vld;
  reg        [50:0]   ways_2_metas_107_tag;
  reg                 ways_2_metas_107_mru;
  reg                 ways_2_metas_108_vld;
  reg        [50:0]   ways_2_metas_108_tag;
  reg                 ways_2_metas_108_mru;
  reg                 ways_2_metas_109_vld;
  reg        [50:0]   ways_2_metas_109_tag;
  reg                 ways_2_metas_109_mru;
  reg                 ways_2_metas_110_vld;
  reg        [50:0]   ways_2_metas_110_tag;
  reg                 ways_2_metas_110_mru;
  reg                 ways_2_metas_111_vld;
  reg        [50:0]   ways_2_metas_111_tag;
  reg                 ways_2_metas_111_mru;
  reg                 ways_2_metas_112_vld;
  reg        [50:0]   ways_2_metas_112_tag;
  reg                 ways_2_metas_112_mru;
  reg                 ways_2_metas_113_vld;
  reg        [50:0]   ways_2_metas_113_tag;
  reg                 ways_2_metas_113_mru;
  reg                 ways_2_metas_114_vld;
  reg        [50:0]   ways_2_metas_114_tag;
  reg                 ways_2_metas_114_mru;
  reg                 ways_2_metas_115_vld;
  reg        [50:0]   ways_2_metas_115_tag;
  reg                 ways_2_metas_115_mru;
  reg                 ways_2_metas_116_vld;
  reg        [50:0]   ways_2_metas_116_tag;
  reg                 ways_2_metas_116_mru;
  reg                 ways_2_metas_117_vld;
  reg        [50:0]   ways_2_metas_117_tag;
  reg                 ways_2_metas_117_mru;
  reg                 ways_2_metas_118_vld;
  reg        [50:0]   ways_2_metas_118_tag;
  reg                 ways_2_metas_118_mru;
  reg                 ways_2_metas_119_vld;
  reg        [50:0]   ways_2_metas_119_tag;
  reg                 ways_2_metas_119_mru;
  reg                 ways_2_metas_120_vld;
  reg        [50:0]   ways_2_metas_120_tag;
  reg                 ways_2_metas_120_mru;
  reg                 ways_2_metas_121_vld;
  reg        [50:0]   ways_2_metas_121_tag;
  reg                 ways_2_metas_121_mru;
  reg                 ways_2_metas_122_vld;
  reg        [50:0]   ways_2_metas_122_tag;
  reg                 ways_2_metas_122_mru;
  reg                 ways_2_metas_123_vld;
  reg        [50:0]   ways_2_metas_123_tag;
  reg                 ways_2_metas_123_mru;
  reg                 ways_2_metas_124_vld;
  reg        [50:0]   ways_2_metas_124_tag;
  reg                 ways_2_metas_124_mru;
  reg                 ways_2_metas_125_vld;
  reg        [50:0]   ways_2_metas_125_tag;
  reg                 ways_2_metas_125_mru;
  reg                 ways_2_metas_126_vld;
  reg        [50:0]   ways_2_metas_126_tag;
  reg                 ways_2_metas_126_mru;
  reg                 ways_2_metas_127_vld;
  reg        [50:0]   ways_2_metas_127_tag;
  reg                 ways_2_metas_127_mru;
  reg                 ways_3_metas_0_vld;
  reg        [50:0]   ways_3_metas_0_tag;
  reg                 ways_3_metas_0_mru;
  reg                 ways_3_metas_1_vld;
  reg        [50:0]   ways_3_metas_1_tag;
  reg                 ways_3_metas_1_mru;
  reg                 ways_3_metas_2_vld;
  reg        [50:0]   ways_3_metas_2_tag;
  reg                 ways_3_metas_2_mru;
  reg                 ways_3_metas_3_vld;
  reg        [50:0]   ways_3_metas_3_tag;
  reg                 ways_3_metas_3_mru;
  reg                 ways_3_metas_4_vld;
  reg        [50:0]   ways_3_metas_4_tag;
  reg                 ways_3_metas_4_mru;
  reg                 ways_3_metas_5_vld;
  reg        [50:0]   ways_3_metas_5_tag;
  reg                 ways_3_metas_5_mru;
  reg                 ways_3_metas_6_vld;
  reg        [50:0]   ways_3_metas_6_tag;
  reg                 ways_3_metas_6_mru;
  reg                 ways_3_metas_7_vld;
  reg        [50:0]   ways_3_metas_7_tag;
  reg                 ways_3_metas_7_mru;
  reg                 ways_3_metas_8_vld;
  reg        [50:0]   ways_3_metas_8_tag;
  reg                 ways_3_metas_8_mru;
  reg                 ways_3_metas_9_vld;
  reg        [50:0]   ways_3_metas_9_tag;
  reg                 ways_3_metas_9_mru;
  reg                 ways_3_metas_10_vld;
  reg        [50:0]   ways_3_metas_10_tag;
  reg                 ways_3_metas_10_mru;
  reg                 ways_3_metas_11_vld;
  reg        [50:0]   ways_3_metas_11_tag;
  reg                 ways_3_metas_11_mru;
  reg                 ways_3_metas_12_vld;
  reg        [50:0]   ways_3_metas_12_tag;
  reg                 ways_3_metas_12_mru;
  reg                 ways_3_metas_13_vld;
  reg        [50:0]   ways_3_metas_13_tag;
  reg                 ways_3_metas_13_mru;
  reg                 ways_3_metas_14_vld;
  reg        [50:0]   ways_3_metas_14_tag;
  reg                 ways_3_metas_14_mru;
  reg                 ways_3_metas_15_vld;
  reg        [50:0]   ways_3_metas_15_tag;
  reg                 ways_3_metas_15_mru;
  reg                 ways_3_metas_16_vld;
  reg        [50:0]   ways_3_metas_16_tag;
  reg                 ways_3_metas_16_mru;
  reg                 ways_3_metas_17_vld;
  reg        [50:0]   ways_3_metas_17_tag;
  reg                 ways_3_metas_17_mru;
  reg                 ways_3_metas_18_vld;
  reg        [50:0]   ways_3_metas_18_tag;
  reg                 ways_3_metas_18_mru;
  reg                 ways_3_metas_19_vld;
  reg        [50:0]   ways_3_metas_19_tag;
  reg                 ways_3_metas_19_mru;
  reg                 ways_3_metas_20_vld;
  reg        [50:0]   ways_3_metas_20_tag;
  reg                 ways_3_metas_20_mru;
  reg                 ways_3_metas_21_vld;
  reg        [50:0]   ways_3_metas_21_tag;
  reg                 ways_3_metas_21_mru;
  reg                 ways_3_metas_22_vld;
  reg        [50:0]   ways_3_metas_22_tag;
  reg                 ways_3_metas_22_mru;
  reg                 ways_3_metas_23_vld;
  reg        [50:0]   ways_3_metas_23_tag;
  reg                 ways_3_metas_23_mru;
  reg                 ways_3_metas_24_vld;
  reg        [50:0]   ways_3_metas_24_tag;
  reg                 ways_3_metas_24_mru;
  reg                 ways_3_metas_25_vld;
  reg        [50:0]   ways_3_metas_25_tag;
  reg                 ways_3_metas_25_mru;
  reg                 ways_3_metas_26_vld;
  reg        [50:0]   ways_3_metas_26_tag;
  reg                 ways_3_metas_26_mru;
  reg                 ways_3_metas_27_vld;
  reg        [50:0]   ways_3_metas_27_tag;
  reg                 ways_3_metas_27_mru;
  reg                 ways_3_metas_28_vld;
  reg        [50:0]   ways_3_metas_28_tag;
  reg                 ways_3_metas_28_mru;
  reg                 ways_3_metas_29_vld;
  reg        [50:0]   ways_3_metas_29_tag;
  reg                 ways_3_metas_29_mru;
  reg                 ways_3_metas_30_vld;
  reg        [50:0]   ways_3_metas_30_tag;
  reg                 ways_3_metas_30_mru;
  reg                 ways_3_metas_31_vld;
  reg        [50:0]   ways_3_metas_31_tag;
  reg                 ways_3_metas_31_mru;
  reg                 ways_3_metas_32_vld;
  reg        [50:0]   ways_3_metas_32_tag;
  reg                 ways_3_metas_32_mru;
  reg                 ways_3_metas_33_vld;
  reg        [50:0]   ways_3_metas_33_tag;
  reg                 ways_3_metas_33_mru;
  reg                 ways_3_metas_34_vld;
  reg        [50:0]   ways_3_metas_34_tag;
  reg                 ways_3_metas_34_mru;
  reg                 ways_3_metas_35_vld;
  reg        [50:0]   ways_3_metas_35_tag;
  reg                 ways_3_metas_35_mru;
  reg                 ways_3_metas_36_vld;
  reg        [50:0]   ways_3_metas_36_tag;
  reg                 ways_3_metas_36_mru;
  reg                 ways_3_metas_37_vld;
  reg        [50:0]   ways_3_metas_37_tag;
  reg                 ways_3_metas_37_mru;
  reg                 ways_3_metas_38_vld;
  reg        [50:0]   ways_3_metas_38_tag;
  reg                 ways_3_metas_38_mru;
  reg                 ways_3_metas_39_vld;
  reg        [50:0]   ways_3_metas_39_tag;
  reg                 ways_3_metas_39_mru;
  reg                 ways_3_metas_40_vld;
  reg        [50:0]   ways_3_metas_40_tag;
  reg                 ways_3_metas_40_mru;
  reg                 ways_3_metas_41_vld;
  reg        [50:0]   ways_3_metas_41_tag;
  reg                 ways_3_metas_41_mru;
  reg                 ways_3_metas_42_vld;
  reg        [50:0]   ways_3_metas_42_tag;
  reg                 ways_3_metas_42_mru;
  reg                 ways_3_metas_43_vld;
  reg        [50:0]   ways_3_metas_43_tag;
  reg                 ways_3_metas_43_mru;
  reg                 ways_3_metas_44_vld;
  reg        [50:0]   ways_3_metas_44_tag;
  reg                 ways_3_metas_44_mru;
  reg                 ways_3_metas_45_vld;
  reg        [50:0]   ways_3_metas_45_tag;
  reg                 ways_3_metas_45_mru;
  reg                 ways_3_metas_46_vld;
  reg        [50:0]   ways_3_metas_46_tag;
  reg                 ways_3_metas_46_mru;
  reg                 ways_3_metas_47_vld;
  reg        [50:0]   ways_3_metas_47_tag;
  reg                 ways_3_metas_47_mru;
  reg                 ways_3_metas_48_vld;
  reg        [50:0]   ways_3_metas_48_tag;
  reg                 ways_3_metas_48_mru;
  reg                 ways_3_metas_49_vld;
  reg        [50:0]   ways_3_metas_49_tag;
  reg                 ways_3_metas_49_mru;
  reg                 ways_3_metas_50_vld;
  reg        [50:0]   ways_3_metas_50_tag;
  reg                 ways_3_metas_50_mru;
  reg                 ways_3_metas_51_vld;
  reg        [50:0]   ways_3_metas_51_tag;
  reg                 ways_3_metas_51_mru;
  reg                 ways_3_metas_52_vld;
  reg        [50:0]   ways_3_metas_52_tag;
  reg                 ways_3_metas_52_mru;
  reg                 ways_3_metas_53_vld;
  reg        [50:0]   ways_3_metas_53_tag;
  reg                 ways_3_metas_53_mru;
  reg                 ways_3_metas_54_vld;
  reg        [50:0]   ways_3_metas_54_tag;
  reg                 ways_3_metas_54_mru;
  reg                 ways_3_metas_55_vld;
  reg        [50:0]   ways_3_metas_55_tag;
  reg                 ways_3_metas_55_mru;
  reg                 ways_3_metas_56_vld;
  reg        [50:0]   ways_3_metas_56_tag;
  reg                 ways_3_metas_56_mru;
  reg                 ways_3_metas_57_vld;
  reg        [50:0]   ways_3_metas_57_tag;
  reg                 ways_3_metas_57_mru;
  reg                 ways_3_metas_58_vld;
  reg        [50:0]   ways_3_metas_58_tag;
  reg                 ways_3_metas_58_mru;
  reg                 ways_3_metas_59_vld;
  reg        [50:0]   ways_3_metas_59_tag;
  reg                 ways_3_metas_59_mru;
  reg                 ways_3_metas_60_vld;
  reg        [50:0]   ways_3_metas_60_tag;
  reg                 ways_3_metas_60_mru;
  reg                 ways_3_metas_61_vld;
  reg        [50:0]   ways_3_metas_61_tag;
  reg                 ways_3_metas_61_mru;
  reg                 ways_3_metas_62_vld;
  reg        [50:0]   ways_3_metas_62_tag;
  reg                 ways_3_metas_62_mru;
  reg                 ways_3_metas_63_vld;
  reg        [50:0]   ways_3_metas_63_tag;
  reg                 ways_3_metas_63_mru;
  reg                 ways_3_metas_64_vld;
  reg        [50:0]   ways_3_metas_64_tag;
  reg                 ways_3_metas_64_mru;
  reg                 ways_3_metas_65_vld;
  reg        [50:0]   ways_3_metas_65_tag;
  reg                 ways_3_metas_65_mru;
  reg                 ways_3_metas_66_vld;
  reg        [50:0]   ways_3_metas_66_tag;
  reg                 ways_3_metas_66_mru;
  reg                 ways_3_metas_67_vld;
  reg        [50:0]   ways_3_metas_67_tag;
  reg                 ways_3_metas_67_mru;
  reg                 ways_3_metas_68_vld;
  reg        [50:0]   ways_3_metas_68_tag;
  reg                 ways_3_metas_68_mru;
  reg                 ways_3_metas_69_vld;
  reg        [50:0]   ways_3_metas_69_tag;
  reg                 ways_3_metas_69_mru;
  reg                 ways_3_metas_70_vld;
  reg        [50:0]   ways_3_metas_70_tag;
  reg                 ways_3_metas_70_mru;
  reg                 ways_3_metas_71_vld;
  reg        [50:0]   ways_3_metas_71_tag;
  reg                 ways_3_metas_71_mru;
  reg                 ways_3_metas_72_vld;
  reg        [50:0]   ways_3_metas_72_tag;
  reg                 ways_3_metas_72_mru;
  reg                 ways_3_metas_73_vld;
  reg        [50:0]   ways_3_metas_73_tag;
  reg                 ways_3_metas_73_mru;
  reg                 ways_3_metas_74_vld;
  reg        [50:0]   ways_3_metas_74_tag;
  reg                 ways_3_metas_74_mru;
  reg                 ways_3_metas_75_vld;
  reg        [50:0]   ways_3_metas_75_tag;
  reg                 ways_3_metas_75_mru;
  reg                 ways_3_metas_76_vld;
  reg        [50:0]   ways_3_metas_76_tag;
  reg                 ways_3_metas_76_mru;
  reg                 ways_3_metas_77_vld;
  reg        [50:0]   ways_3_metas_77_tag;
  reg                 ways_3_metas_77_mru;
  reg                 ways_3_metas_78_vld;
  reg        [50:0]   ways_3_metas_78_tag;
  reg                 ways_3_metas_78_mru;
  reg                 ways_3_metas_79_vld;
  reg        [50:0]   ways_3_metas_79_tag;
  reg                 ways_3_metas_79_mru;
  reg                 ways_3_metas_80_vld;
  reg        [50:0]   ways_3_metas_80_tag;
  reg                 ways_3_metas_80_mru;
  reg                 ways_3_metas_81_vld;
  reg        [50:0]   ways_3_metas_81_tag;
  reg                 ways_3_metas_81_mru;
  reg                 ways_3_metas_82_vld;
  reg        [50:0]   ways_3_metas_82_tag;
  reg                 ways_3_metas_82_mru;
  reg                 ways_3_metas_83_vld;
  reg        [50:0]   ways_3_metas_83_tag;
  reg                 ways_3_metas_83_mru;
  reg                 ways_3_metas_84_vld;
  reg        [50:0]   ways_3_metas_84_tag;
  reg                 ways_3_metas_84_mru;
  reg                 ways_3_metas_85_vld;
  reg        [50:0]   ways_3_metas_85_tag;
  reg                 ways_3_metas_85_mru;
  reg                 ways_3_metas_86_vld;
  reg        [50:0]   ways_3_metas_86_tag;
  reg                 ways_3_metas_86_mru;
  reg                 ways_3_metas_87_vld;
  reg        [50:0]   ways_3_metas_87_tag;
  reg                 ways_3_metas_87_mru;
  reg                 ways_3_metas_88_vld;
  reg        [50:0]   ways_3_metas_88_tag;
  reg                 ways_3_metas_88_mru;
  reg                 ways_3_metas_89_vld;
  reg        [50:0]   ways_3_metas_89_tag;
  reg                 ways_3_metas_89_mru;
  reg                 ways_3_metas_90_vld;
  reg        [50:0]   ways_3_metas_90_tag;
  reg                 ways_3_metas_90_mru;
  reg                 ways_3_metas_91_vld;
  reg        [50:0]   ways_3_metas_91_tag;
  reg                 ways_3_metas_91_mru;
  reg                 ways_3_metas_92_vld;
  reg        [50:0]   ways_3_metas_92_tag;
  reg                 ways_3_metas_92_mru;
  reg                 ways_3_metas_93_vld;
  reg        [50:0]   ways_3_metas_93_tag;
  reg                 ways_3_metas_93_mru;
  reg                 ways_3_metas_94_vld;
  reg        [50:0]   ways_3_metas_94_tag;
  reg                 ways_3_metas_94_mru;
  reg                 ways_3_metas_95_vld;
  reg        [50:0]   ways_3_metas_95_tag;
  reg                 ways_3_metas_95_mru;
  reg                 ways_3_metas_96_vld;
  reg        [50:0]   ways_3_metas_96_tag;
  reg                 ways_3_metas_96_mru;
  reg                 ways_3_metas_97_vld;
  reg        [50:0]   ways_3_metas_97_tag;
  reg                 ways_3_metas_97_mru;
  reg                 ways_3_metas_98_vld;
  reg        [50:0]   ways_3_metas_98_tag;
  reg                 ways_3_metas_98_mru;
  reg                 ways_3_metas_99_vld;
  reg        [50:0]   ways_3_metas_99_tag;
  reg                 ways_3_metas_99_mru;
  reg                 ways_3_metas_100_vld;
  reg        [50:0]   ways_3_metas_100_tag;
  reg                 ways_3_metas_100_mru;
  reg                 ways_3_metas_101_vld;
  reg        [50:0]   ways_3_metas_101_tag;
  reg                 ways_3_metas_101_mru;
  reg                 ways_3_metas_102_vld;
  reg        [50:0]   ways_3_metas_102_tag;
  reg                 ways_3_metas_102_mru;
  reg                 ways_3_metas_103_vld;
  reg        [50:0]   ways_3_metas_103_tag;
  reg                 ways_3_metas_103_mru;
  reg                 ways_3_metas_104_vld;
  reg        [50:0]   ways_3_metas_104_tag;
  reg                 ways_3_metas_104_mru;
  reg                 ways_3_metas_105_vld;
  reg        [50:0]   ways_3_metas_105_tag;
  reg                 ways_3_metas_105_mru;
  reg                 ways_3_metas_106_vld;
  reg        [50:0]   ways_3_metas_106_tag;
  reg                 ways_3_metas_106_mru;
  reg                 ways_3_metas_107_vld;
  reg        [50:0]   ways_3_metas_107_tag;
  reg                 ways_3_metas_107_mru;
  reg                 ways_3_metas_108_vld;
  reg        [50:0]   ways_3_metas_108_tag;
  reg                 ways_3_metas_108_mru;
  reg                 ways_3_metas_109_vld;
  reg        [50:0]   ways_3_metas_109_tag;
  reg                 ways_3_metas_109_mru;
  reg                 ways_3_metas_110_vld;
  reg        [50:0]   ways_3_metas_110_tag;
  reg                 ways_3_metas_110_mru;
  reg                 ways_3_metas_111_vld;
  reg        [50:0]   ways_3_metas_111_tag;
  reg                 ways_3_metas_111_mru;
  reg                 ways_3_metas_112_vld;
  reg        [50:0]   ways_3_metas_112_tag;
  reg                 ways_3_metas_112_mru;
  reg                 ways_3_metas_113_vld;
  reg        [50:0]   ways_3_metas_113_tag;
  reg                 ways_3_metas_113_mru;
  reg                 ways_3_metas_114_vld;
  reg        [50:0]   ways_3_metas_114_tag;
  reg                 ways_3_metas_114_mru;
  reg                 ways_3_metas_115_vld;
  reg        [50:0]   ways_3_metas_115_tag;
  reg                 ways_3_metas_115_mru;
  reg                 ways_3_metas_116_vld;
  reg        [50:0]   ways_3_metas_116_tag;
  reg                 ways_3_metas_116_mru;
  reg                 ways_3_metas_117_vld;
  reg        [50:0]   ways_3_metas_117_tag;
  reg                 ways_3_metas_117_mru;
  reg                 ways_3_metas_118_vld;
  reg        [50:0]   ways_3_metas_118_tag;
  reg                 ways_3_metas_118_mru;
  reg                 ways_3_metas_119_vld;
  reg        [50:0]   ways_3_metas_119_tag;
  reg                 ways_3_metas_119_mru;
  reg                 ways_3_metas_120_vld;
  reg        [50:0]   ways_3_metas_120_tag;
  reg                 ways_3_metas_120_mru;
  reg                 ways_3_metas_121_vld;
  reg        [50:0]   ways_3_metas_121_tag;
  reg                 ways_3_metas_121_mru;
  reg                 ways_3_metas_122_vld;
  reg        [50:0]   ways_3_metas_122_tag;
  reg                 ways_3_metas_122_mru;
  reg                 ways_3_metas_123_vld;
  reg        [50:0]   ways_3_metas_123_tag;
  reg                 ways_3_metas_123_mru;
  reg                 ways_3_metas_124_vld;
  reg        [50:0]   ways_3_metas_124_tag;
  reg                 ways_3_metas_124_mru;
  reg                 ways_3_metas_125_vld;
  reg        [50:0]   ways_3_metas_125_tag;
  reg                 ways_3_metas_125_mru;
  reg                 ways_3_metas_126_vld;
  reg        [50:0]   ways_3_metas_126_tag;
  reg                 ways_3_metas_126_mru;
  reg                 ways_3_metas_127_vld;
  reg        [50:0]   ways_3_metas_127_tag;
  reg                 ways_3_metas_127_mru;
  wire       [50:0]   cache_tag_0;
  wire       [50:0]   cache_tag_1;
  wire       [50:0]   cache_tag_2;
  wire       [50:0]   cache_tag_3;
  wire                cache_hit_0;
  wire                cache_hit_1;
  wire                cache_hit_2;
  wire                cache_hit_3;
  wire                cache_invld_d1_0;
  wire                cache_invld_d1_1;
  wire                cache_invld_d1_2;
  wire                cache_invld_d1_3;
  wire                cache_victim_0;
  wire                cache_victim_1;
  wire                cache_victim_2;
  wire                cache_victim_3;
  wire                cache_mru_0;
  wire                cache_mru_1;
  wire                cache_mru_2;
  wire                cache_mru_3;
  wire                cache_lru_d1_0;
  wire                cache_lru_d1_1;
  wire                cache_lru_d1_2;
  wire                cache_lru_d1_3;
  wire       [1:0]    hit_id;
  reg        [1:0]    hit_id_d1;
  wire       [1:0]    evict_id;
  wire       [1:0]    invld_id;
  wire       [1:0]    victim_id;
  wire                mru_full;
  wire                cpu_cmd_fire;
  wire                is_hit;
  reg                 is_hit_d1;
  wire                cpu_cmd_fire_1;
  wire                is_miss;
  wire                is_diff;
  reg                 flush_busy;
  reg                 flush_cnt_willIncrement;
  reg                 flush_cnt_willClear;
  reg        [6:0]    flush_cnt_valueNext;
  reg        [6:0]    flush_cnt_value;
  wire                flush_cnt_willOverflowIfInc;
  wire                flush_cnt_willOverflow;
  wire                flush_done;
  wire                cache_hit_gnt_0;
  wire                cache_hit_gnt_1;
  wire                cache_hit_gnt_2;
  wire                cache_hit_gnt_3;
  wire                cache_victim_gnt_0;
  wire                cache_victim_gnt_1;
  wire                cache_victim_gnt_2;
  wire                cache_victim_gnt_3;
  wire                cache_invld_gnt_0;
  wire                cache_invld_gnt_1;
  wire                cache_invld_gnt_2;
  wire                cache_invld_gnt_3;
  reg        [1:0]    evict_id_miss;
  wire       [50:0]   cpu_tag;
  wire       [6:0]    cpu_set;
  wire       [6:0]    cpu_bank_addr;
  wire       [3:0]    cpu_bank_index;
  wire                cpu_cmd_fire_2;
  reg        [63:0]   cpu_addr_d1;
  wire       [6:0]    cpu_set_d1;
  wire       [50:0]   cpu_tag_d1;
  wire       [6:0]    cpu_bank_addr_d1;
  wire       [3:0]    cpu_bank_index_d1;
  reg                 cpu_cmd_ready_1;
  wire       [511:0]  sram_banks_data_0;
  wire       [511:0]  sram_banks_data_1;
  wire       [511:0]  sram_banks_data_2;
  wire       [511:0]  sram_banks_data_3;
  wire                sram_banks_valid_0;
  wire                sram_banks_valid_1;
  wire                sram_banks_valid_2;
  wire                sram_banks_valid_3;
  reg                 next_level_cmd_valid_1;
  reg                 next_level_data_cnt_willIncrement;
  reg                 next_level_data_cnt_willClear;
  reg        [2:0]    next_level_data_cnt_valueNext;
  reg        [2:0]    next_level_data_cnt_value;
  wire                next_level_data_cnt_willOverflowIfInc;
  wire                next_level_data_cnt_willOverflow;
  wire       [6:0]    next_level_bank_addr;
  reg                 next_level_done;
  wire                next_level_cmd_fire;
  wire                when_ICache_l142;
  wire       [3:0]    _zz_cache_hit_gnt_0;
  wire       [3:0]    _zz_cache_hit_gnt_0_1;
  wire       [7:0]    _zz_cache_hit_gnt_0_2;
  wire       [7:0]    _zz_cache_hit_gnt_0_3;
  wire       [3:0]    _zz_cache_hit_gnt_0_4;
  wire       [3:0]    _zz_cache_invld_gnt_0;
  wire       [3:0]    _zz_cache_invld_gnt_0_1;
  wire       [7:0]    _zz_cache_invld_gnt_0_2;
  wire       [7:0]    _zz_cache_invld_gnt_0_3;
  wire       [3:0]    _zz_cache_invld_gnt_0_4;
  wire       [3:0]    _zz_cache_victim_gnt_0;
  wire       [3:0]    _zz_cache_victim_gnt_0_1;
  wire       [7:0]    _zz_cache_victim_gnt_0_2;
  wire       [7:0]    _zz_cache_victim_gnt_0_3;
  wire       [3:0]    _zz_cache_victim_gnt_0_4;
  wire                _zz_hit_id;
  wire                _zz_hit_id_1;
  wire                _zz_invld_id;
  wire                _zz_invld_id_1;
  wire                _zz_victim_id;
  wire                _zz_victim_id_1;
  wire       [127:0]  _zz_1;
  wire                _zz_2;
  wire                _zz_3;
  wire                _zz_4;
  wire                _zz_5;
  wire                _zz_6;
  wire                _zz_7;
  wire                _zz_8;
  wire                _zz_9;
  wire                _zz_10;
  wire                _zz_11;
  wire                _zz_12;
  wire                _zz_13;
  wire                _zz_14;
  wire                _zz_15;
  wire                _zz_16;
  wire                _zz_17;
  wire                _zz_18;
  wire                _zz_19;
  wire                _zz_20;
  wire                _zz_21;
  wire                _zz_22;
  wire                _zz_23;
  wire                _zz_24;
  wire                _zz_25;
  wire                _zz_26;
  wire                _zz_27;
  wire                _zz_28;
  wire                _zz_29;
  wire                _zz_30;
  wire                _zz_31;
  wire                _zz_32;
  wire                _zz_33;
  wire                _zz_34;
  wire                _zz_35;
  wire                _zz_36;
  wire                _zz_37;
  wire                _zz_38;
  wire                _zz_39;
  wire                _zz_40;
  wire                _zz_41;
  wire                _zz_42;
  wire                _zz_43;
  wire                _zz_44;
  wire                _zz_45;
  wire                _zz_46;
  wire                _zz_47;
  wire                _zz_48;
  wire                _zz_49;
  wire                _zz_50;
  wire                _zz_51;
  wire                _zz_52;
  wire                _zz_53;
  wire                _zz_54;
  wire                _zz_55;
  wire                _zz_56;
  wire                _zz_57;
  wire                _zz_58;
  wire                _zz_59;
  wire                _zz_60;
  wire                _zz_61;
  wire                _zz_62;
  wire                _zz_63;
  wire                _zz_64;
  wire                _zz_65;
  wire                _zz_66;
  wire                _zz_67;
  wire                _zz_68;
  wire                _zz_69;
  wire                _zz_70;
  wire                _zz_71;
  wire                _zz_72;
  wire                _zz_73;
  wire                _zz_74;
  wire                _zz_75;
  wire                _zz_76;
  wire                _zz_77;
  wire                _zz_78;
  wire                _zz_79;
  wire                _zz_80;
  wire                _zz_81;
  wire                _zz_82;
  wire                _zz_83;
  wire                _zz_84;
  wire                _zz_85;
  wire                _zz_86;
  wire                _zz_87;
  wire                _zz_88;
  wire                _zz_89;
  wire                _zz_90;
  wire                _zz_91;
  wire                _zz_92;
  wire                _zz_93;
  wire                _zz_94;
  wire                _zz_95;
  wire                _zz_96;
  wire                _zz_97;
  wire                _zz_98;
  wire                _zz_99;
  wire                _zz_100;
  wire                _zz_101;
  wire                _zz_102;
  wire                _zz_103;
  wire                _zz_104;
  wire                _zz_105;
  wire                _zz_106;
  wire                _zz_107;
  wire                _zz_108;
  wire                _zz_109;
  wire                _zz_110;
  wire                _zz_111;
  wire                _zz_112;
  wire                _zz_113;
  wire                _zz_114;
  wire                _zz_115;
  wire                _zz_116;
  wire                _zz_117;
  wire                _zz_118;
  wire                _zz_119;
  wire                _zz_120;
  wire                _zz_121;
  wire                _zz_122;
  wire                _zz_123;
  wire                _zz_124;
  wire                _zz_125;
  wire                _zz_126;
  wire                _zz_127;
  wire                _zz_128;
  wire                _zz_129;
  wire       [127:0]  _zz_130;
  wire                _zz_131;
  wire                _zz_132;
  wire                _zz_133;
  wire                _zz_134;
  wire                _zz_135;
  wire                _zz_136;
  wire                _zz_137;
  wire                _zz_138;
  wire                _zz_139;
  wire                _zz_140;
  wire                _zz_141;
  wire                _zz_142;
  wire                _zz_143;
  wire                _zz_144;
  wire                _zz_145;
  wire                _zz_146;
  wire                _zz_147;
  wire                _zz_148;
  wire                _zz_149;
  wire                _zz_150;
  wire                _zz_151;
  wire                _zz_152;
  wire                _zz_153;
  wire                _zz_154;
  wire                _zz_155;
  wire                _zz_156;
  wire                _zz_157;
  wire                _zz_158;
  wire                _zz_159;
  wire                _zz_160;
  wire                _zz_161;
  wire                _zz_162;
  wire                _zz_163;
  wire                _zz_164;
  wire                _zz_165;
  wire                _zz_166;
  wire                _zz_167;
  wire                _zz_168;
  wire                _zz_169;
  wire                _zz_170;
  wire                _zz_171;
  wire                _zz_172;
  wire                _zz_173;
  wire                _zz_174;
  wire                _zz_175;
  wire                _zz_176;
  wire                _zz_177;
  wire                _zz_178;
  wire                _zz_179;
  wire                _zz_180;
  wire                _zz_181;
  wire                _zz_182;
  wire                _zz_183;
  wire                _zz_184;
  wire                _zz_185;
  wire                _zz_186;
  wire                _zz_187;
  wire                _zz_188;
  wire                _zz_189;
  wire                _zz_190;
  wire                _zz_191;
  wire                _zz_192;
  wire                _zz_193;
  wire                _zz_194;
  wire                _zz_195;
  wire                _zz_196;
  wire                _zz_197;
  wire                _zz_198;
  wire                _zz_199;
  wire                _zz_200;
  wire                _zz_201;
  wire                _zz_202;
  wire                _zz_203;
  wire                _zz_204;
  wire                _zz_205;
  wire                _zz_206;
  wire                _zz_207;
  wire                _zz_208;
  wire                _zz_209;
  wire                _zz_210;
  wire                _zz_211;
  wire                _zz_212;
  wire                _zz_213;
  wire                _zz_214;
  wire                _zz_215;
  wire                _zz_216;
  wire                _zz_217;
  wire                _zz_218;
  wire                _zz_219;
  wire                _zz_220;
  wire                _zz_221;
  wire                _zz_222;
  wire                _zz_223;
  wire                _zz_224;
  wire                _zz_225;
  wire                _zz_226;
  wire                _zz_227;
  wire                _zz_228;
  wire                _zz_229;
  wire                _zz_230;
  wire                _zz_231;
  wire                _zz_232;
  wire                _zz_233;
  wire                _zz_234;
  wire                _zz_235;
  wire                _zz_236;
  wire                _zz_237;
  wire                _zz_238;
  wire                _zz_239;
  wire                _zz_240;
  wire                _zz_241;
  wire                _zz_242;
  wire                _zz_243;
  wire                _zz_244;
  wire                _zz_245;
  wire                _zz_246;
  wire                _zz_247;
  wire                _zz_248;
  wire                _zz_249;
  wire                _zz_250;
  wire                _zz_251;
  wire                _zz_252;
  wire                _zz_253;
  wire                _zz_254;
  wire                _zz_255;
  wire                _zz_256;
  wire                _zz_257;
  wire                _zz_258;
  wire                when_ICache_l174;
  reg        [15:0]   _zz_sram_0_ports_cmd_payload_wen;
  wire                when_ICache_l181;
  wire                when_ICache_l188;
  wire       [127:0]  _zz_259;
  wire                _zz_260;
  wire                _zz_261;
  wire                _zz_262;
  wire                _zz_263;
  wire                _zz_264;
  wire                _zz_265;
  wire                _zz_266;
  wire                _zz_267;
  wire                _zz_268;
  wire                _zz_269;
  wire                _zz_270;
  wire                _zz_271;
  wire                _zz_272;
  wire                _zz_273;
  wire                _zz_274;
  wire                _zz_275;
  wire                _zz_276;
  wire                _zz_277;
  wire                _zz_278;
  wire                _zz_279;
  wire                _zz_280;
  wire                _zz_281;
  wire                _zz_282;
  wire                _zz_283;
  wire                _zz_284;
  wire                _zz_285;
  wire                _zz_286;
  wire                _zz_287;
  wire                _zz_288;
  wire                _zz_289;
  wire                _zz_290;
  wire                _zz_291;
  wire                _zz_292;
  wire                _zz_293;
  wire                _zz_294;
  wire                _zz_295;
  wire                _zz_296;
  wire                _zz_297;
  wire                _zz_298;
  wire                _zz_299;
  wire                _zz_300;
  wire                _zz_301;
  wire                _zz_302;
  wire                _zz_303;
  wire                _zz_304;
  wire                _zz_305;
  wire                _zz_306;
  wire                _zz_307;
  wire                _zz_308;
  wire                _zz_309;
  wire                _zz_310;
  wire                _zz_311;
  wire                _zz_312;
  wire                _zz_313;
  wire                _zz_314;
  wire                _zz_315;
  wire                _zz_316;
  wire                _zz_317;
  wire                _zz_318;
  wire                _zz_319;
  wire                _zz_320;
  wire                _zz_321;
  wire                _zz_322;
  wire                _zz_323;
  wire                _zz_324;
  wire                _zz_325;
  wire                _zz_326;
  wire                _zz_327;
  wire                _zz_328;
  wire                _zz_329;
  wire                _zz_330;
  wire                _zz_331;
  wire                _zz_332;
  wire                _zz_333;
  wire                _zz_334;
  wire                _zz_335;
  wire                _zz_336;
  wire                _zz_337;
  wire                _zz_338;
  wire                _zz_339;
  wire                _zz_340;
  wire                _zz_341;
  wire                _zz_342;
  wire                _zz_343;
  wire                _zz_344;
  wire                _zz_345;
  wire                _zz_346;
  wire                _zz_347;
  wire                _zz_348;
  wire                _zz_349;
  wire                _zz_350;
  wire                _zz_351;
  wire                _zz_352;
  wire                _zz_353;
  wire                _zz_354;
  wire                _zz_355;
  wire                _zz_356;
  wire                _zz_357;
  wire                _zz_358;
  wire                _zz_359;
  wire                _zz_360;
  wire                _zz_361;
  wire                _zz_362;
  wire                _zz_363;
  wire                _zz_364;
  wire                _zz_365;
  wire                _zz_366;
  wire                _zz_367;
  wire                _zz_368;
  wire                _zz_369;
  wire                _zz_370;
  wire                _zz_371;
  wire                _zz_372;
  wire                _zz_373;
  wire                _zz_374;
  wire                _zz_375;
  wire                _zz_376;
  wire                _zz_377;
  wire                _zz_378;
  wire                _zz_379;
  wire                _zz_380;
  wire                _zz_381;
  wire                _zz_382;
  wire                _zz_383;
  wire                _zz_384;
  wire                _zz_385;
  wire                _zz_386;
  wire                _zz_387;
  wire                when_ICache_l210;
  wire                when_ICache_l217;
  wire                when_ICache_l220;
  wire                when_ICache_l225;
  wire                when_ICache_l230;
  wire                when_ICache_l233;
  wire       [127:0]  _zz_388;
  wire                _zz_389;
  wire                _zz_390;
  wire                _zz_391;
  wire                _zz_392;
  wire                _zz_393;
  wire                _zz_394;
  wire                _zz_395;
  wire                _zz_396;
  wire                _zz_397;
  wire                _zz_398;
  wire                _zz_399;
  wire                _zz_400;
  wire                _zz_401;
  wire                _zz_402;
  wire                _zz_403;
  wire                _zz_404;
  wire                _zz_405;
  wire                _zz_406;
  wire                _zz_407;
  wire                _zz_408;
  wire                _zz_409;
  wire                _zz_410;
  wire                _zz_411;
  wire                _zz_412;
  wire                _zz_413;
  wire                _zz_414;
  wire                _zz_415;
  wire                _zz_416;
  wire                _zz_417;
  wire                _zz_418;
  wire                _zz_419;
  wire                _zz_420;
  wire                _zz_421;
  wire                _zz_422;
  wire                _zz_423;
  wire                _zz_424;
  wire                _zz_425;
  wire                _zz_426;
  wire                _zz_427;
  wire                _zz_428;
  wire                _zz_429;
  wire                _zz_430;
  wire                _zz_431;
  wire                _zz_432;
  wire                _zz_433;
  wire                _zz_434;
  wire                _zz_435;
  wire                _zz_436;
  wire                _zz_437;
  wire                _zz_438;
  wire                _zz_439;
  wire                _zz_440;
  wire                _zz_441;
  wire                _zz_442;
  wire                _zz_443;
  wire                _zz_444;
  wire                _zz_445;
  wire                _zz_446;
  wire                _zz_447;
  wire                _zz_448;
  wire                _zz_449;
  wire                _zz_450;
  wire                _zz_451;
  wire                _zz_452;
  wire                _zz_453;
  wire                _zz_454;
  wire                _zz_455;
  wire                _zz_456;
  wire                _zz_457;
  wire                _zz_458;
  wire                _zz_459;
  wire                _zz_460;
  wire                _zz_461;
  wire                _zz_462;
  wire                _zz_463;
  wire                _zz_464;
  wire                _zz_465;
  wire                _zz_466;
  wire                _zz_467;
  wire                _zz_468;
  wire                _zz_469;
  wire                _zz_470;
  wire                _zz_471;
  wire                _zz_472;
  wire                _zz_473;
  wire                _zz_474;
  wire                _zz_475;
  wire                _zz_476;
  wire                _zz_477;
  wire                _zz_478;
  wire                _zz_479;
  wire                _zz_480;
  wire                _zz_481;
  wire                _zz_482;
  wire                _zz_483;
  wire                _zz_484;
  wire                _zz_485;
  wire                _zz_486;
  wire                _zz_487;
  wire                _zz_488;
  wire                _zz_489;
  wire                _zz_490;
  wire                _zz_491;
  wire                _zz_492;
  wire                _zz_493;
  wire                _zz_494;
  wire                _zz_495;
  wire                _zz_496;
  wire                _zz_497;
  wire                _zz_498;
  wire                _zz_499;
  wire                _zz_500;
  wire                _zz_501;
  wire                _zz_502;
  wire                _zz_503;
  wire                _zz_504;
  wire                _zz_505;
  wire                _zz_506;
  wire                _zz_507;
  wire                _zz_508;
  wire                _zz_509;
  wire                _zz_510;
  wire                _zz_511;
  wire                _zz_512;
  wire                _zz_513;
  wire                _zz_514;
  wire                _zz_515;
  wire                _zz_516;
  wire       [127:0]  _zz_517;
  wire                _zz_518;
  wire                _zz_519;
  wire                _zz_520;
  wire                _zz_521;
  wire                _zz_522;
  wire                _zz_523;
  wire                _zz_524;
  wire                _zz_525;
  wire                _zz_526;
  wire                _zz_527;
  wire                _zz_528;
  wire                _zz_529;
  wire                _zz_530;
  wire                _zz_531;
  wire                _zz_532;
  wire                _zz_533;
  wire                _zz_534;
  wire                _zz_535;
  wire                _zz_536;
  wire                _zz_537;
  wire                _zz_538;
  wire                _zz_539;
  wire                _zz_540;
  wire                _zz_541;
  wire                _zz_542;
  wire                _zz_543;
  wire                _zz_544;
  wire                _zz_545;
  wire                _zz_546;
  wire                _zz_547;
  wire                _zz_548;
  wire                _zz_549;
  wire                _zz_550;
  wire                _zz_551;
  wire                _zz_552;
  wire                _zz_553;
  wire                _zz_554;
  wire                _zz_555;
  wire                _zz_556;
  wire                _zz_557;
  wire                _zz_558;
  wire                _zz_559;
  wire                _zz_560;
  wire                _zz_561;
  wire                _zz_562;
  wire                _zz_563;
  wire                _zz_564;
  wire                _zz_565;
  wire                _zz_566;
  wire                _zz_567;
  wire                _zz_568;
  wire                _zz_569;
  wire                _zz_570;
  wire                _zz_571;
  wire                _zz_572;
  wire                _zz_573;
  wire                _zz_574;
  wire                _zz_575;
  wire                _zz_576;
  wire                _zz_577;
  wire                _zz_578;
  wire                _zz_579;
  wire                _zz_580;
  wire                _zz_581;
  wire                _zz_582;
  wire                _zz_583;
  wire                _zz_584;
  wire                _zz_585;
  wire                _zz_586;
  wire                _zz_587;
  wire                _zz_588;
  wire                _zz_589;
  wire                _zz_590;
  wire                _zz_591;
  wire                _zz_592;
  wire                _zz_593;
  wire                _zz_594;
  wire                _zz_595;
  wire                _zz_596;
  wire                _zz_597;
  wire                _zz_598;
  wire                _zz_599;
  wire                _zz_600;
  wire                _zz_601;
  wire                _zz_602;
  wire                _zz_603;
  wire                _zz_604;
  wire                _zz_605;
  wire                _zz_606;
  wire                _zz_607;
  wire                _zz_608;
  wire                _zz_609;
  wire                _zz_610;
  wire                _zz_611;
  wire                _zz_612;
  wire                _zz_613;
  wire                _zz_614;
  wire                _zz_615;
  wire                _zz_616;
  wire                _zz_617;
  wire                _zz_618;
  wire                _zz_619;
  wire                _zz_620;
  wire                _zz_621;
  wire                _zz_622;
  wire                _zz_623;
  wire                _zz_624;
  wire                _zz_625;
  wire                _zz_626;
  wire                _zz_627;
  wire                _zz_628;
  wire                _zz_629;
  wire                _zz_630;
  wire                _zz_631;
  wire                _zz_632;
  wire                _zz_633;
  wire                _zz_634;
  wire                _zz_635;
  wire                _zz_636;
  wire                _zz_637;
  wire                _zz_638;
  wire                _zz_639;
  wire                _zz_640;
  wire                _zz_641;
  wire                _zz_642;
  wire                _zz_643;
  wire                _zz_644;
  wire                _zz_645;
  wire                when_ICache_l174_1;
  reg        [15:0]   _zz_sram_1_ports_cmd_payload_wen;
  wire                when_ICache_l181_1;
  wire                when_ICache_l188_1;
  wire       [127:0]  _zz_646;
  wire                _zz_647;
  wire                _zz_648;
  wire                _zz_649;
  wire                _zz_650;
  wire                _zz_651;
  wire                _zz_652;
  wire                _zz_653;
  wire                _zz_654;
  wire                _zz_655;
  wire                _zz_656;
  wire                _zz_657;
  wire                _zz_658;
  wire                _zz_659;
  wire                _zz_660;
  wire                _zz_661;
  wire                _zz_662;
  wire                _zz_663;
  wire                _zz_664;
  wire                _zz_665;
  wire                _zz_666;
  wire                _zz_667;
  wire                _zz_668;
  wire                _zz_669;
  wire                _zz_670;
  wire                _zz_671;
  wire                _zz_672;
  wire                _zz_673;
  wire                _zz_674;
  wire                _zz_675;
  wire                _zz_676;
  wire                _zz_677;
  wire                _zz_678;
  wire                _zz_679;
  wire                _zz_680;
  wire                _zz_681;
  wire                _zz_682;
  wire                _zz_683;
  wire                _zz_684;
  wire                _zz_685;
  wire                _zz_686;
  wire                _zz_687;
  wire                _zz_688;
  wire                _zz_689;
  wire                _zz_690;
  wire                _zz_691;
  wire                _zz_692;
  wire                _zz_693;
  wire                _zz_694;
  wire                _zz_695;
  wire                _zz_696;
  wire                _zz_697;
  wire                _zz_698;
  wire                _zz_699;
  wire                _zz_700;
  wire                _zz_701;
  wire                _zz_702;
  wire                _zz_703;
  wire                _zz_704;
  wire                _zz_705;
  wire                _zz_706;
  wire                _zz_707;
  wire                _zz_708;
  wire                _zz_709;
  wire                _zz_710;
  wire                _zz_711;
  wire                _zz_712;
  wire                _zz_713;
  wire                _zz_714;
  wire                _zz_715;
  wire                _zz_716;
  wire                _zz_717;
  wire                _zz_718;
  wire                _zz_719;
  wire                _zz_720;
  wire                _zz_721;
  wire                _zz_722;
  wire                _zz_723;
  wire                _zz_724;
  wire                _zz_725;
  wire                _zz_726;
  wire                _zz_727;
  wire                _zz_728;
  wire                _zz_729;
  wire                _zz_730;
  wire                _zz_731;
  wire                _zz_732;
  wire                _zz_733;
  wire                _zz_734;
  wire                _zz_735;
  wire                _zz_736;
  wire                _zz_737;
  wire                _zz_738;
  wire                _zz_739;
  wire                _zz_740;
  wire                _zz_741;
  wire                _zz_742;
  wire                _zz_743;
  wire                _zz_744;
  wire                _zz_745;
  wire                _zz_746;
  wire                _zz_747;
  wire                _zz_748;
  wire                _zz_749;
  wire                _zz_750;
  wire                _zz_751;
  wire                _zz_752;
  wire                _zz_753;
  wire                _zz_754;
  wire                _zz_755;
  wire                _zz_756;
  wire                _zz_757;
  wire                _zz_758;
  wire                _zz_759;
  wire                _zz_760;
  wire                _zz_761;
  wire                _zz_762;
  wire                _zz_763;
  wire                _zz_764;
  wire                _zz_765;
  wire                _zz_766;
  wire                _zz_767;
  wire                _zz_768;
  wire                _zz_769;
  wire                _zz_770;
  wire                _zz_771;
  wire                _zz_772;
  wire                _zz_773;
  wire                _zz_774;
  wire                when_ICache_l210_1;
  wire                when_ICache_l217_1;
  wire                when_ICache_l220_1;
  wire                when_ICache_l225_1;
  wire                when_ICache_l230_1;
  wire                when_ICache_l233_1;
  wire       [127:0]  _zz_775;
  wire                _zz_776;
  wire                _zz_777;
  wire                _zz_778;
  wire                _zz_779;
  wire                _zz_780;
  wire                _zz_781;
  wire                _zz_782;
  wire                _zz_783;
  wire                _zz_784;
  wire                _zz_785;
  wire                _zz_786;
  wire                _zz_787;
  wire                _zz_788;
  wire                _zz_789;
  wire                _zz_790;
  wire                _zz_791;
  wire                _zz_792;
  wire                _zz_793;
  wire                _zz_794;
  wire                _zz_795;
  wire                _zz_796;
  wire                _zz_797;
  wire                _zz_798;
  wire                _zz_799;
  wire                _zz_800;
  wire                _zz_801;
  wire                _zz_802;
  wire                _zz_803;
  wire                _zz_804;
  wire                _zz_805;
  wire                _zz_806;
  wire                _zz_807;
  wire                _zz_808;
  wire                _zz_809;
  wire                _zz_810;
  wire                _zz_811;
  wire                _zz_812;
  wire                _zz_813;
  wire                _zz_814;
  wire                _zz_815;
  wire                _zz_816;
  wire                _zz_817;
  wire                _zz_818;
  wire                _zz_819;
  wire                _zz_820;
  wire                _zz_821;
  wire                _zz_822;
  wire                _zz_823;
  wire                _zz_824;
  wire                _zz_825;
  wire                _zz_826;
  wire                _zz_827;
  wire                _zz_828;
  wire                _zz_829;
  wire                _zz_830;
  wire                _zz_831;
  wire                _zz_832;
  wire                _zz_833;
  wire                _zz_834;
  wire                _zz_835;
  wire                _zz_836;
  wire                _zz_837;
  wire                _zz_838;
  wire                _zz_839;
  wire                _zz_840;
  wire                _zz_841;
  wire                _zz_842;
  wire                _zz_843;
  wire                _zz_844;
  wire                _zz_845;
  wire                _zz_846;
  wire                _zz_847;
  wire                _zz_848;
  wire                _zz_849;
  wire                _zz_850;
  wire                _zz_851;
  wire                _zz_852;
  wire                _zz_853;
  wire                _zz_854;
  wire                _zz_855;
  wire                _zz_856;
  wire                _zz_857;
  wire                _zz_858;
  wire                _zz_859;
  wire                _zz_860;
  wire                _zz_861;
  wire                _zz_862;
  wire                _zz_863;
  wire                _zz_864;
  wire                _zz_865;
  wire                _zz_866;
  wire                _zz_867;
  wire                _zz_868;
  wire                _zz_869;
  wire                _zz_870;
  wire                _zz_871;
  wire                _zz_872;
  wire                _zz_873;
  wire                _zz_874;
  wire                _zz_875;
  wire                _zz_876;
  wire                _zz_877;
  wire                _zz_878;
  wire                _zz_879;
  wire                _zz_880;
  wire                _zz_881;
  wire                _zz_882;
  wire                _zz_883;
  wire                _zz_884;
  wire                _zz_885;
  wire                _zz_886;
  wire                _zz_887;
  wire                _zz_888;
  wire                _zz_889;
  wire                _zz_890;
  wire                _zz_891;
  wire                _zz_892;
  wire                _zz_893;
  wire                _zz_894;
  wire                _zz_895;
  wire                _zz_896;
  wire                _zz_897;
  wire                _zz_898;
  wire                _zz_899;
  wire                _zz_900;
  wire                _zz_901;
  wire                _zz_902;
  wire                _zz_903;
  wire       [127:0]  _zz_904;
  wire                _zz_905;
  wire                _zz_906;
  wire                _zz_907;
  wire                _zz_908;
  wire                _zz_909;
  wire                _zz_910;
  wire                _zz_911;
  wire                _zz_912;
  wire                _zz_913;
  wire                _zz_914;
  wire                _zz_915;
  wire                _zz_916;
  wire                _zz_917;
  wire                _zz_918;
  wire                _zz_919;
  wire                _zz_920;
  wire                _zz_921;
  wire                _zz_922;
  wire                _zz_923;
  wire                _zz_924;
  wire                _zz_925;
  wire                _zz_926;
  wire                _zz_927;
  wire                _zz_928;
  wire                _zz_929;
  wire                _zz_930;
  wire                _zz_931;
  wire                _zz_932;
  wire                _zz_933;
  wire                _zz_934;
  wire                _zz_935;
  wire                _zz_936;
  wire                _zz_937;
  wire                _zz_938;
  wire                _zz_939;
  wire                _zz_940;
  wire                _zz_941;
  wire                _zz_942;
  wire                _zz_943;
  wire                _zz_944;
  wire                _zz_945;
  wire                _zz_946;
  wire                _zz_947;
  wire                _zz_948;
  wire                _zz_949;
  wire                _zz_950;
  wire                _zz_951;
  wire                _zz_952;
  wire                _zz_953;
  wire                _zz_954;
  wire                _zz_955;
  wire                _zz_956;
  wire                _zz_957;
  wire                _zz_958;
  wire                _zz_959;
  wire                _zz_960;
  wire                _zz_961;
  wire                _zz_962;
  wire                _zz_963;
  wire                _zz_964;
  wire                _zz_965;
  wire                _zz_966;
  wire                _zz_967;
  wire                _zz_968;
  wire                _zz_969;
  wire                _zz_970;
  wire                _zz_971;
  wire                _zz_972;
  wire                _zz_973;
  wire                _zz_974;
  wire                _zz_975;
  wire                _zz_976;
  wire                _zz_977;
  wire                _zz_978;
  wire                _zz_979;
  wire                _zz_980;
  wire                _zz_981;
  wire                _zz_982;
  wire                _zz_983;
  wire                _zz_984;
  wire                _zz_985;
  wire                _zz_986;
  wire                _zz_987;
  wire                _zz_988;
  wire                _zz_989;
  wire                _zz_990;
  wire                _zz_991;
  wire                _zz_992;
  wire                _zz_993;
  wire                _zz_994;
  wire                _zz_995;
  wire                _zz_996;
  wire                _zz_997;
  wire                _zz_998;
  wire                _zz_999;
  wire                _zz_1000;
  wire                _zz_1001;
  wire                _zz_1002;
  wire                _zz_1003;
  wire                _zz_1004;
  wire                _zz_1005;
  wire                _zz_1006;
  wire                _zz_1007;
  wire                _zz_1008;
  wire                _zz_1009;
  wire                _zz_1010;
  wire                _zz_1011;
  wire                _zz_1012;
  wire                _zz_1013;
  wire                _zz_1014;
  wire                _zz_1015;
  wire                _zz_1016;
  wire                _zz_1017;
  wire                _zz_1018;
  wire                _zz_1019;
  wire                _zz_1020;
  wire                _zz_1021;
  wire                _zz_1022;
  wire                _zz_1023;
  wire                _zz_1024;
  wire                _zz_1025;
  wire                _zz_1026;
  wire                _zz_1027;
  wire                _zz_1028;
  wire                _zz_1029;
  wire                _zz_1030;
  wire                _zz_1031;
  wire                _zz_1032;
  wire                when_ICache_l174_2;
  reg        [15:0]   _zz_sram_2_ports_cmd_payload_wen;
  wire                when_ICache_l181_2;
  wire                when_ICache_l188_2;
  wire       [127:0]  _zz_1033;
  wire                _zz_1034;
  wire                _zz_1035;
  wire                _zz_1036;
  wire                _zz_1037;
  wire                _zz_1038;
  wire                _zz_1039;
  wire                _zz_1040;
  wire                _zz_1041;
  wire                _zz_1042;
  wire                _zz_1043;
  wire                _zz_1044;
  wire                _zz_1045;
  wire                _zz_1046;
  wire                _zz_1047;
  wire                _zz_1048;
  wire                _zz_1049;
  wire                _zz_1050;
  wire                _zz_1051;
  wire                _zz_1052;
  wire                _zz_1053;
  wire                _zz_1054;
  wire                _zz_1055;
  wire                _zz_1056;
  wire                _zz_1057;
  wire                _zz_1058;
  wire                _zz_1059;
  wire                _zz_1060;
  wire                _zz_1061;
  wire                _zz_1062;
  wire                _zz_1063;
  wire                _zz_1064;
  wire                _zz_1065;
  wire                _zz_1066;
  wire                _zz_1067;
  wire                _zz_1068;
  wire                _zz_1069;
  wire                _zz_1070;
  wire                _zz_1071;
  wire                _zz_1072;
  wire                _zz_1073;
  wire                _zz_1074;
  wire                _zz_1075;
  wire                _zz_1076;
  wire                _zz_1077;
  wire                _zz_1078;
  wire                _zz_1079;
  wire                _zz_1080;
  wire                _zz_1081;
  wire                _zz_1082;
  wire                _zz_1083;
  wire                _zz_1084;
  wire                _zz_1085;
  wire                _zz_1086;
  wire                _zz_1087;
  wire                _zz_1088;
  wire                _zz_1089;
  wire                _zz_1090;
  wire                _zz_1091;
  wire                _zz_1092;
  wire                _zz_1093;
  wire                _zz_1094;
  wire                _zz_1095;
  wire                _zz_1096;
  wire                _zz_1097;
  wire                _zz_1098;
  wire                _zz_1099;
  wire                _zz_1100;
  wire                _zz_1101;
  wire                _zz_1102;
  wire                _zz_1103;
  wire                _zz_1104;
  wire                _zz_1105;
  wire                _zz_1106;
  wire                _zz_1107;
  wire                _zz_1108;
  wire                _zz_1109;
  wire                _zz_1110;
  wire                _zz_1111;
  wire                _zz_1112;
  wire                _zz_1113;
  wire                _zz_1114;
  wire                _zz_1115;
  wire                _zz_1116;
  wire                _zz_1117;
  wire                _zz_1118;
  wire                _zz_1119;
  wire                _zz_1120;
  wire                _zz_1121;
  wire                _zz_1122;
  wire                _zz_1123;
  wire                _zz_1124;
  wire                _zz_1125;
  wire                _zz_1126;
  wire                _zz_1127;
  wire                _zz_1128;
  wire                _zz_1129;
  wire                _zz_1130;
  wire                _zz_1131;
  wire                _zz_1132;
  wire                _zz_1133;
  wire                _zz_1134;
  wire                _zz_1135;
  wire                _zz_1136;
  wire                _zz_1137;
  wire                _zz_1138;
  wire                _zz_1139;
  wire                _zz_1140;
  wire                _zz_1141;
  wire                _zz_1142;
  wire                _zz_1143;
  wire                _zz_1144;
  wire                _zz_1145;
  wire                _zz_1146;
  wire                _zz_1147;
  wire                _zz_1148;
  wire                _zz_1149;
  wire                _zz_1150;
  wire                _zz_1151;
  wire                _zz_1152;
  wire                _zz_1153;
  wire                _zz_1154;
  wire                _zz_1155;
  wire                _zz_1156;
  wire                _zz_1157;
  wire                _zz_1158;
  wire                _zz_1159;
  wire                _zz_1160;
  wire                _zz_1161;
  wire                when_ICache_l210_2;
  wire                when_ICache_l217_2;
  wire                when_ICache_l220_2;
  wire                when_ICache_l225_2;
  wire                when_ICache_l230_2;
  wire                when_ICache_l233_2;
  wire       [127:0]  _zz_1162;
  wire                _zz_1163;
  wire                _zz_1164;
  wire                _zz_1165;
  wire                _zz_1166;
  wire                _zz_1167;
  wire                _zz_1168;
  wire                _zz_1169;
  wire                _zz_1170;
  wire                _zz_1171;
  wire                _zz_1172;
  wire                _zz_1173;
  wire                _zz_1174;
  wire                _zz_1175;
  wire                _zz_1176;
  wire                _zz_1177;
  wire                _zz_1178;
  wire                _zz_1179;
  wire                _zz_1180;
  wire                _zz_1181;
  wire                _zz_1182;
  wire                _zz_1183;
  wire                _zz_1184;
  wire                _zz_1185;
  wire                _zz_1186;
  wire                _zz_1187;
  wire                _zz_1188;
  wire                _zz_1189;
  wire                _zz_1190;
  wire                _zz_1191;
  wire                _zz_1192;
  wire                _zz_1193;
  wire                _zz_1194;
  wire                _zz_1195;
  wire                _zz_1196;
  wire                _zz_1197;
  wire                _zz_1198;
  wire                _zz_1199;
  wire                _zz_1200;
  wire                _zz_1201;
  wire                _zz_1202;
  wire                _zz_1203;
  wire                _zz_1204;
  wire                _zz_1205;
  wire                _zz_1206;
  wire                _zz_1207;
  wire                _zz_1208;
  wire                _zz_1209;
  wire                _zz_1210;
  wire                _zz_1211;
  wire                _zz_1212;
  wire                _zz_1213;
  wire                _zz_1214;
  wire                _zz_1215;
  wire                _zz_1216;
  wire                _zz_1217;
  wire                _zz_1218;
  wire                _zz_1219;
  wire                _zz_1220;
  wire                _zz_1221;
  wire                _zz_1222;
  wire                _zz_1223;
  wire                _zz_1224;
  wire                _zz_1225;
  wire                _zz_1226;
  wire                _zz_1227;
  wire                _zz_1228;
  wire                _zz_1229;
  wire                _zz_1230;
  wire                _zz_1231;
  wire                _zz_1232;
  wire                _zz_1233;
  wire                _zz_1234;
  wire                _zz_1235;
  wire                _zz_1236;
  wire                _zz_1237;
  wire                _zz_1238;
  wire                _zz_1239;
  wire                _zz_1240;
  wire                _zz_1241;
  wire                _zz_1242;
  wire                _zz_1243;
  wire                _zz_1244;
  wire                _zz_1245;
  wire                _zz_1246;
  wire                _zz_1247;
  wire                _zz_1248;
  wire                _zz_1249;
  wire                _zz_1250;
  wire                _zz_1251;
  wire                _zz_1252;
  wire                _zz_1253;
  wire                _zz_1254;
  wire                _zz_1255;
  wire                _zz_1256;
  wire                _zz_1257;
  wire                _zz_1258;
  wire                _zz_1259;
  wire                _zz_1260;
  wire                _zz_1261;
  wire                _zz_1262;
  wire                _zz_1263;
  wire                _zz_1264;
  wire                _zz_1265;
  wire                _zz_1266;
  wire                _zz_1267;
  wire                _zz_1268;
  wire                _zz_1269;
  wire                _zz_1270;
  wire                _zz_1271;
  wire                _zz_1272;
  wire                _zz_1273;
  wire                _zz_1274;
  wire                _zz_1275;
  wire                _zz_1276;
  wire                _zz_1277;
  wire                _zz_1278;
  wire                _zz_1279;
  wire                _zz_1280;
  wire                _zz_1281;
  wire                _zz_1282;
  wire                _zz_1283;
  wire                _zz_1284;
  wire                _zz_1285;
  wire                _zz_1286;
  wire                _zz_1287;
  wire                _zz_1288;
  wire                _zz_1289;
  wire                _zz_1290;
  wire       [127:0]  _zz_1291;
  wire                _zz_1292;
  wire                _zz_1293;
  wire                _zz_1294;
  wire                _zz_1295;
  wire                _zz_1296;
  wire                _zz_1297;
  wire                _zz_1298;
  wire                _zz_1299;
  wire                _zz_1300;
  wire                _zz_1301;
  wire                _zz_1302;
  wire                _zz_1303;
  wire                _zz_1304;
  wire                _zz_1305;
  wire                _zz_1306;
  wire                _zz_1307;
  wire                _zz_1308;
  wire                _zz_1309;
  wire                _zz_1310;
  wire                _zz_1311;
  wire                _zz_1312;
  wire                _zz_1313;
  wire                _zz_1314;
  wire                _zz_1315;
  wire                _zz_1316;
  wire                _zz_1317;
  wire                _zz_1318;
  wire                _zz_1319;
  wire                _zz_1320;
  wire                _zz_1321;
  wire                _zz_1322;
  wire                _zz_1323;
  wire                _zz_1324;
  wire                _zz_1325;
  wire                _zz_1326;
  wire                _zz_1327;
  wire                _zz_1328;
  wire                _zz_1329;
  wire                _zz_1330;
  wire                _zz_1331;
  wire                _zz_1332;
  wire                _zz_1333;
  wire                _zz_1334;
  wire                _zz_1335;
  wire                _zz_1336;
  wire                _zz_1337;
  wire                _zz_1338;
  wire                _zz_1339;
  wire                _zz_1340;
  wire                _zz_1341;
  wire                _zz_1342;
  wire                _zz_1343;
  wire                _zz_1344;
  wire                _zz_1345;
  wire                _zz_1346;
  wire                _zz_1347;
  wire                _zz_1348;
  wire                _zz_1349;
  wire                _zz_1350;
  wire                _zz_1351;
  wire                _zz_1352;
  wire                _zz_1353;
  wire                _zz_1354;
  wire                _zz_1355;
  wire                _zz_1356;
  wire                _zz_1357;
  wire                _zz_1358;
  wire                _zz_1359;
  wire                _zz_1360;
  wire                _zz_1361;
  wire                _zz_1362;
  wire                _zz_1363;
  wire                _zz_1364;
  wire                _zz_1365;
  wire                _zz_1366;
  wire                _zz_1367;
  wire                _zz_1368;
  wire                _zz_1369;
  wire                _zz_1370;
  wire                _zz_1371;
  wire                _zz_1372;
  wire                _zz_1373;
  wire                _zz_1374;
  wire                _zz_1375;
  wire                _zz_1376;
  wire                _zz_1377;
  wire                _zz_1378;
  wire                _zz_1379;
  wire                _zz_1380;
  wire                _zz_1381;
  wire                _zz_1382;
  wire                _zz_1383;
  wire                _zz_1384;
  wire                _zz_1385;
  wire                _zz_1386;
  wire                _zz_1387;
  wire                _zz_1388;
  wire                _zz_1389;
  wire                _zz_1390;
  wire                _zz_1391;
  wire                _zz_1392;
  wire                _zz_1393;
  wire                _zz_1394;
  wire                _zz_1395;
  wire                _zz_1396;
  wire                _zz_1397;
  wire                _zz_1398;
  wire                _zz_1399;
  wire                _zz_1400;
  wire                _zz_1401;
  wire                _zz_1402;
  wire                _zz_1403;
  wire                _zz_1404;
  wire                _zz_1405;
  wire                _zz_1406;
  wire                _zz_1407;
  wire                _zz_1408;
  wire                _zz_1409;
  wire                _zz_1410;
  wire                _zz_1411;
  wire                _zz_1412;
  wire                _zz_1413;
  wire                _zz_1414;
  wire                _zz_1415;
  wire                _zz_1416;
  wire                _zz_1417;
  wire                _zz_1418;
  wire                _zz_1419;
  wire                when_ICache_l174_3;
  reg        [15:0]   _zz_sram_3_ports_cmd_payload_wen;
  wire                when_ICache_l181_3;
  wire                when_ICache_l188_3;
  wire       [127:0]  _zz_1420;
  wire                _zz_1421;
  wire                _zz_1422;
  wire                _zz_1423;
  wire                _zz_1424;
  wire                _zz_1425;
  wire                _zz_1426;
  wire                _zz_1427;
  wire                _zz_1428;
  wire                _zz_1429;
  wire                _zz_1430;
  wire                _zz_1431;
  wire                _zz_1432;
  wire                _zz_1433;
  wire                _zz_1434;
  wire                _zz_1435;
  wire                _zz_1436;
  wire                _zz_1437;
  wire                _zz_1438;
  wire                _zz_1439;
  wire                _zz_1440;
  wire                _zz_1441;
  wire                _zz_1442;
  wire                _zz_1443;
  wire                _zz_1444;
  wire                _zz_1445;
  wire                _zz_1446;
  wire                _zz_1447;
  wire                _zz_1448;
  wire                _zz_1449;
  wire                _zz_1450;
  wire                _zz_1451;
  wire                _zz_1452;
  wire                _zz_1453;
  wire                _zz_1454;
  wire                _zz_1455;
  wire                _zz_1456;
  wire                _zz_1457;
  wire                _zz_1458;
  wire                _zz_1459;
  wire                _zz_1460;
  wire                _zz_1461;
  wire                _zz_1462;
  wire                _zz_1463;
  wire                _zz_1464;
  wire                _zz_1465;
  wire                _zz_1466;
  wire                _zz_1467;
  wire                _zz_1468;
  wire                _zz_1469;
  wire                _zz_1470;
  wire                _zz_1471;
  wire                _zz_1472;
  wire                _zz_1473;
  wire                _zz_1474;
  wire                _zz_1475;
  wire                _zz_1476;
  wire                _zz_1477;
  wire                _zz_1478;
  wire                _zz_1479;
  wire                _zz_1480;
  wire                _zz_1481;
  wire                _zz_1482;
  wire                _zz_1483;
  wire                _zz_1484;
  wire                _zz_1485;
  wire                _zz_1486;
  wire                _zz_1487;
  wire                _zz_1488;
  wire                _zz_1489;
  wire                _zz_1490;
  wire                _zz_1491;
  wire                _zz_1492;
  wire                _zz_1493;
  wire                _zz_1494;
  wire                _zz_1495;
  wire                _zz_1496;
  wire                _zz_1497;
  wire                _zz_1498;
  wire                _zz_1499;
  wire                _zz_1500;
  wire                _zz_1501;
  wire                _zz_1502;
  wire                _zz_1503;
  wire                _zz_1504;
  wire                _zz_1505;
  wire                _zz_1506;
  wire                _zz_1507;
  wire                _zz_1508;
  wire                _zz_1509;
  wire                _zz_1510;
  wire                _zz_1511;
  wire                _zz_1512;
  wire                _zz_1513;
  wire                _zz_1514;
  wire                _zz_1515;
  wire                _zz_1516;
  wire                _zz_1517;
  wire                _zz_1518;
  wire                _zz_1519;
  wire                _zz_1520;
  wire                _zz_1521;
  wire                _zz_1522;
  wire                _zz_1523;
  wire                _zz_1524;
  wire                _zz_1525;
  wire                _zz_1526;
  wire                _zz_1527;
  wire                _zz_1528;
  wire                _zz_1529;
  wire                _zz_1530;
  wire                _zz_1531;
  wire                _zz_1532;
  wire                _zz_1533;
  wire                _zz_1534;
  wire                _zz_1535;
  wire                _zz_1536;
  wire                _zz_1537;
  wire                _zz_1538;
  wire                _zz_1539;
  wire                _zz_1540;
  wire                _zz_1541;
  wire                _zz_1542;
  wire                _zz_1543;
  wire                _zz_1544;
  wire                _zz_1545;
  wire                _zz_1546;
  wire                _zz_1547;
  wire                _zz_1548;
  wire                when_ICache_l210_3;
  wire                when_ICache_l217_3;
  wire                when_ICache_l220_3;
  wire                when_ICache_l225_3;
  wire                when_ICache_l230_3;
  wire                when_ICache_l233_3;
  wire       [511:0]  _zz_cpu_rsp_payload_data;
  wire       [511:0]  _zz_cpu_rsp_payload_data_1;
  function [15:0] zz__zz_sram_0_ports_cmd_payload_wen(input dummy);
    begin
      zz__zz_sram_0_ports_cmd_payload_wen = 16'h0;
      zz__zz_sram_0_ports_cmd_payload_wen[1] = 1'b1;
      zz__zz_sram_0_ports_cmd_payload_wen[0] = 1'b1;
    end
  endfunction
  wire [15:0] _zz_1549;
  function [15:0] zz__zz_sram_1_ports_cmd_payload_wen(input dummy);
    begin
      zz__zz_sram_1_ports_cmd_payload_wen = 16'h0;
      zz__zz_sram_1_ports_cmd_payload_wen[1] = 1'b1;
      zz__zz_sram_1_ports_cmd_payload_wen[0] = 1'b1;
    end
  endfunction
  wire [15:0] _zz_1550;
  function [15:0] zz__zz_sram_2_ports_cmd_payload_wen(input dummy);
    begin
      zz__zz_sram_2_ports_cmd_payload_wen = 16'h0;
      zz__zz_sram_2_ports_cmd_payload_wen[1] = 1'b1;
      zz__zz_sram_2_ports_cmd_payload_wen[0] = 1'b1;
    end
  endfunction
  wire [15:0] _zz_1551;
  function [15:0] zz__zz_sram_3_ports_cmd_payload_wen(input dummy);
    begin
      zz__zz_sram_3_ports_cmd_payload_wen = 16'h0;
      zz__zz_sram_3_ports_cmd_payload_wen[1] = 1'b1;
      zz__zz_sram_3_ports_cmd_payload_wen[0] = 1'b1;
    end
  endfunction
  wire [15:0] _zz_1552;

  assign _zz_flush_cnt_valueNext_1 = flush_cnt_willIncrement;
  assign _zz_flush_cnt_valueNext = {6'd0, _zz_flush_cnt_valueNext_1};
  assign _zz_next_level_data_cnt_valueNext_1 = next_level_data_cnt_willIncrement;
  assign _zz_next_level_data_cnt_valueNext = {2'd0, _zz_next_level_data_cnt_valueNext_1};
  assign _zz__zz_cache_hit_gnt_0_3 = (_zz_cache_hit_gnt_0_2 - _zz__zz_cache_hit_gnt_0_3_1);
  assign _zz__zz_cache_hit_gnt_0_3_2 = {_zz_cache_hit_gnt_0[3],{_zz_cache_hit_gnt_0[2],{_zz_cache_hit_gnt_0[1],_zz_cache_hit_gnt_0[0]}}};
  assign _zz__zz_cache_hit_gnt_0_3_1 = {4'd0, _zz__zz_cache_hit_gnt_0_3_2};
  assign _zz__zz_cache_invld_gnt_0_3 = (_zz_cache_invld_gnt_0_2 - _zz__zz_cache_invld_gnt_0_3_1);
  assign _zz__zz_cache_invld_gnt_0_3_2 = {_zz_cache_invld_gnt_0[3],{_zz_cache_invld_gnt_0[2],{_zz_cache_invld_gnt_0[1],_zz_cache_invld_gnt_0[0]}}};
  assign _zz__zz_cache_invld_gnt_0_3_1 = {4'd0, _zz__zz_cache_invld_gnt_0_3_2};
  assign _zz__zz_cache_victim_gnt_0_3 = (_zz_cache_victim_gnt_0_2 - _zz__zz_cache_victim_gnt_0_3_1);
  assign _zz__zz_cache_victim_gnt_0_3_2 = {_zz_cache_victim_gnt_0[3],{_zz_cache_victim_gnt_0[2],{_zz_cache_victim_gnt_0[1],_zz_cache_victim_gnt_0[0]}}};
  assign _zz__zz_cache_victim_gnt_0_3_1 = {4'd0, _zz__zz_cache_victim_gnt_0_3_2};
  assign _zz_sram_0_ports_cmd_payload_wen_1 = (next_level_data_cnt_value * 2'b10);
  assign _zz_sram_0_ports_cmd_payload_wdata = (next_level_data_cnt_value * 7'h40);
  assign _zz_sram_0_ports_cmd_payload_wstrb = (_zz_sram_0_ports_cmd_payload_wstrb_1 / 4'b1000);
  assign _zz_sram_0_ports_cmd_payload_wstrb_1 = (next_level_data_cnt_value * 7'h40);
  assign _zz_sram_1_ports_cmd_payload_wen_1 = (next_level_data_cnt_value * 2'b10);
  assign _zz_sram_1_ports_cmd_payload_wdata = (next_level_data_cnt_value * 7'h40);
  assign _zz_sram_1_ports_cmd_payload_wstrb = (_zz_sram_1_ports_cmd_payload_wstrb_1 / 4'b1000);
  assign _zz_sram_1_ports_cmd_payload_wstrb_1 = (next_level_data_cnt_value * 7'h40);
  assign _zz_sram_2_ports_cmd_payload_wen_1 = (next_level_data_cnt_value * 2'b10);
  assign _zz_sram_2_ports_cmd_payload_wdata = (next_level_data_cnt_value * 7'h40);
  assign _zz_sram_2_ports_cmd_payload_wstrb = (_zz_sram_2_ports_cmd_payload_wstrb_1 / 4'b1000);
  assign _zz_sram_2_ports_cmd_payload_wstrb_1 = (next_level_data_cnt_value * 7'h40);
  assign _zz_sram_3_ports_cmd_payload_wen_1 = (next_level_data_cnt_value * 2'b10);
  assign _zz_sram_3_ports_cmd_payload_wdata = (next_level_data_cnt_value * 7'h40);
  assign _zz_sram_3_ports_cmd_payload_wstrb = (_zz_sram_3_ports_cmd_payload_wstrb_1 / 4'b1000);
  assign _zz_sram_3_ports_cmd_payload_wstrb_1 = (next_level_data_cnt_value * 7'h40);
  always @(*) begin
    case(cpu_set)
      7'b0000000 : begin
        _zz_cache_tag_0 = ways_0_metas_0_tag;
        _zz_cache_hit_0 = ways_0_metas_0_vld;
        _zz_cache_mru_0 = ways_0_metas_0_mru;
        _zz_cache_tag_1 = ways_1_metas_0_tag;
        _zz_cache_hit_1 = ways_1_metas_0_vld;
        _zz_cache_mru_1 = ways_1_metas_0_mru;
        _zz_cache_tag_2 = ways_2_metas_0_tag;
        _zz_cache_hit_2 = ways_2_metas_0_vld;
        _zz_cache_mru_2 = ways_2_metas_0_mru;
        _zz_cache_tag_3 = ways_3_metas_0_tag;
        _zz_cache_hit_3 = ways_3_metas_0_vld;
        _zz_cache_mru_3 = ways_3_metas_0_mru;
      end
      7'b0000001 : begin
        _zz_cache_tag_0 = ways_0_metas_1_tag;
        _zz_cache_hit_0 = ways_0_metas_1_vld;
        _zz_cache_mru_0 = ways_0_metas_1_mru;
        _zz_cache_tag_1 = ways_1_metas_1_tag;
        _zz_cache_hit_1 = ways_1_metas_1_vld;
        _zz_cache_mru_1 = ways_1_metas_1_mru;
        _zz_cache_tag_2 = ways_2_metas_1_tag;
        _zz_cache_hit_2 = ways_2_metas_1_vld;
        _zz_cache_mru_2 = ways_2_metas_1_mru;
        _zz_cache_tag_3 = ways_3_metas_1_tag;
        _zz_cache_hit_3 = ways_3_metas_1_vld;
        _zz_cache_mru_3 = ways_3_metas_1_mru;
      end
      7'b0000010 : begin
        _zz_cache_tag_0 = ways_0_metas_2_tag;
        _zz_cache_hit_0 = ways_0_metas_2_vld;
        _zz_cache_mru_0 = ways_0_metas_2_mru;
        _zz_cache_tag_1 = ways_1_metas_2_tag;
        _zz_cache_hit_1 = ways_1_metas_2_vld;
        _zz_cache_mru_1 = ways_1_metas_2_mru;
        _zz_cache_tag_2 = ways_2_metas_2_tag;
        _zz_cache_hit_2 = ways_2_metas_2_vld;
        _zz_cache_mru_2 = ways_2_metas_2_mru;
        _zz_cache_tag_3 = ways_3_metas_2_tag;
        _zz_cache_hit_3 = ways_3_metas_2_vld;
        _zz_cache_mru_3 = ways_3_metas_2_mru;
      end
      7'b0000011 : begin
        _zz_cache_tag_0 = ways_0_metas_3_tag;
        _zz_cache_hit_0 = ways_0_metas_3_vld;
        _zz_cache_mru_0 = ways_0_metas_3_mru;
        _zz_cache_tag_1 = ways_1_metas_3_tag;
        _zz_cache_hit_1 = ways_1_metas_3_vld;
        _zz_cache_mru_1 = ways_1_metas_3_mru;
        _zz_cache_tag_2 = ways_2_metas_3_tag;
        _zz_cache_hit_2 = ways_2_metas_3_vld;
        _zz_cache_mru_2 = ways_2_metas_3_mru;
        _zz_cache_tag_3 = ways_3_metas_3_tag;
        _zz_cache_hit_3 = ways_3_metas_3_vld;
        _zz_cache_mru_3 = ways_3_metas_3_mru;
      end
      7'b0000100 : begin
        _zz_cache_tag_0 = ways_0_metas_4_tag;
        _zz_cache_hit_0 = ways_0_metas_4_vld;
        _zz_cache_mru_0 = ways_0_metas_4_mru;
        _zz_cache_tag_1 = ways_1_metas_4_tag;
        _zz_cache_hit_1 = ways_1_metas_4_vld;
        _zz_cache_mru_1 = ways_1_metas_4_mru;
        _zz_cache_tag_2 = ways_2_metas_4_tag;
        _zz_cache_hit_2 = ways_2_metas_4_vld;
        _zz_cache_mru_2 = ways_2_metas_4_mru;
        _zz_cache_tag_3 = ways_3_metas_4_tag;
        _zz_cache_hit_3 = ways_3_metas_4_vld;
        _zz_cache_mru_3 = ways_3_metas_4_mru;
      end
      7'b0000101 : begin
        _zz_cache_tag_0 = ways_0_metas_5_tag;
        _zz_cache_hit_0 = ways_0_metas_5_vld;
        _zz_cache_mru_0 = ways_0_metas_5_mru;
        _zz_cache_tag_1 = ways_1_metas_5_tag;
        _zz_cache_hit_1 = ways_1_metas_5_vld;
        _zz_cache_mru_1 = ways_1_metas_5_mru;
        _zz_cache_tag_2 = ways_2_metas_5_tag;
        _zz_cache_hit_2 = ways_2_metas_5_vld;
        _zz_cache_mru_2 = ways_2_metas_5_mru;
        _zz_cache_tag_3 = ways_3_metas_5_tag;
        _zz_cache_hit_3 = ways_3_metas_5_vld;
        _zz_cache_mru_3 = ways_3_metas_5_mru;
      end
      7'b0000110 : begin
        _zz_cache_tag_0 = ways_0_metas_6_tag;
        _zz_cache_hit_0 = ways_0_metas_6_vld;
        _zz_cache_mru_0 = ways_0_metas_6_mru;
        _zz_cache_tag_1 = ways_1_metas_6_tag;
        _zz_cache_hit_1 = ways_1_metas_6_vld;
        _zz_cache_mru_1 = ways_1_metas_6_mru;
        _zz_cache_tag_2 = ways_2_metas_6_tag;
        _zz_cache_hit_2 = ways_2_metas_6_vld;
        _zz_cache_mru_2 = ways_2_metas_6_mru;
        _zz_cache_tag_3 = ways_3_metas_6_tag;
        _zz_cache_hit_3 = ways_3_metas_6_vld;
        _zz_cache_mru_3 = ways_3_metas_6_mru;
      end
      7'b0000111 : begin
        _zz_cache_tag_0 = ways_0_metas_7_tag;
        _zz_cache_hit_0 = ways_0_metas_7_vld;
        _zz_cache_mru_0 = ways_0_metas_7_mru;
        _zz_cache_tag_1 = ways_1_metas_7_tag;
        _zz_cache_hit_1 = ways_1_metas_7_vld;
        _zz_cache_mru_1 = ways_1_metas_7_mru;
        _zz_cache_tag_2 = ways_2_metas_7_tag;
        _zz_cache_hit_2 = ways_2_metas_7_vld;
        _zz_cache_mru_2 = ways_2_metas_7_mru;
        _zz_cache_tag_3 = ways_3_metas_7_tag;
        _zz_cache_hit_3 = ways_3_metas_7_vld;
        _zz_cache_mru_3 = ways_3_metas_7_mru;
      end
      7'b0001000 : begin
        _zz_cache_tag_0 = ways_0_metas_8_tag;
        _zz_cache_hit_0 = ways_0_metas_8_vld;
        _zz_cache_mru_0 = ways_0_metas_8_mru;
        _zz_cache_tag_1 = ways_1_metas_8_tag;
        _zz_cache_hit_1 = ways_1_metas_8_vld;
        _zz_cache_mru_1 = ways_1_metas_8_mru;
        _zz_cache_tag_2 = ways_2_metas_8_tag;
        _zz_cache_hit_2 = ways_2_metas_8_vld;
        _zz_cache_mru_2 = ways_2_metas_8_mru;
        _zz_cache_tag_3 = ways_3_metas_8_tag;
        _zz_cache_hit_3 = ways_3_metas_8_vld;
        _zz_cache_mru_3 = ways_3_metas_8_mru;
      end
      7'b0001001 : begin
        _zz_cache_tag_0 = ways_0_metas_9_tag;
        _zz_cache_hit_0 = ways_0_metas_9_vld;
        _zz_cache_mru_0 = ways_0_metas_9_mru;
        _zz_cache_tag_1 = ways_1_metas_9_tag;
        _zz_cache_hit_1 = ways_1_metas_9_vld;
        _zz_cache_mru_1 = ways_1_metas_9_mru;
        _zz_cache_tag_2 = ways_2_metas_9_tag;
        _zz_cache_hit_2 = ways_2_metas_9_vld;
        _zz_cache_mru_2 = ways_2_metas_9_mru;
        _zz_cache_tag_3 = ways_3_metas_9_tag;
        _zz_cache_hit_3 = ways_3_metas_9_vld;
        _zz_cache_mru_3 = ways_3_metas_9_mru;
      end
      7'b0001010 : begin
        _zz_cache_tag_0 = ways_0_metas_10_tag;
        _zz_cache_hit_0 = ways_0_metas_10_vld;
        _zz_cache_mru_0 = ways_0_metas_10_mru;
        _zz_cache_tag_1 = ways_1_metas_10_tag;
        _zz_cache_hit_1 = ways_1_metas_10_vld;
        _zz_cache_mru_1 = ways_1_metas_10_mru;
        _zz_cache_tag_2 = ways_2_metas_10_tag;
        _zz_cache_hit_2 = ways_2_metas_10_vld;
        _zz_cache_mru_2 = ways_2_metas_10_mru;
        _zz_cache_tag_3 = ways_3_metas_10_tag;
        _zz_cache_hit_3 = ways_3_metas_10_vld;
        _zz_cache_mru_3 = ways_3_metas_10_mru;
      end
      7'b0001011 : begin
        _zz_cache_tag_0 = ways_0_metas_11_tag;
        _zz_cache_hit_0 = ways_0_metas_11_vld;
        _zz_cache_mru_0 = ways_0_metas_11_mru;
        _zz_cache_tag_1 = ways_1_metas_11_tag;
        _zz_cache_hit_1 = ways_1_metas_11_vld;
        _zz_cache_mru_1 = ways_1_metas_11_mru;
        _zz_cache_tag_2 = ways_2_metas_11_tag;
        _zz_cache_hit_2 = ways_2_metas_11_vld;
        _zz_cache_mru_2 = ways_2_metas_11_mru;
        _zz_cache_tag_3 = ways_3_metas_11_tag;
        _zz_cache_hit_3 = ways_3_metas_11_vld;
        _zz_cache_mru_3 = ways_3_metas_11_mru;
      end
      7'b0001100 : begin
        _zz_cache_tag_0 = ways_0_metas_12_tag;
        _zz_cache_hit_0 = ways_0_metas_12_vld;
        _zz_cache_mru_0 = ways_0_metas_12_mru;
        _zz_cache_tag_1 = ways_1_metas_12_tag;
        _zz_cache_hit_1 = ways_1_metas_12_vld;
        _zz_cache_mru_1 = ways_1_metas_12_mru;
        _zz_cache_tag_2 = ways_2_metas_12_tag;
        _zz_cache_hit_2 = ways_2_metas_12_vld;
        _zz_cache_mru_2 = ways_2_metas_12_mru;
        _zz_cache_tag_3 = ways_3_metas_12_tag;
        _zz_cache_hit_3 = ways_3_metas_12_vld;
        _zz_cache_mru_3 = ways_3_metas_12_mru;
      end
      7'b0001101 : begin
        _zz_cache_tag_0 = ways_0_metas_13_tag;
        _zz_cache_hit_0 = ways_0_metas_13_vld;
        _zz_cache_mru_0 = ways_0_metas_13_mru;
        _zz_cache_tag_1 = ways_1_metas_13_tag;
        _zz_cache_hit_1 = ways_1_metas_13_vld;
        _zz_cache_mru_1 = ways_1_metas_13_mru;
        _zz_cache_tag_2 = ways_2_metas_13_tag;
        _zz_cache_hit_2 = ways_2_metas_13_vld;
        _zz_cache_mru_2 = ways_2_metas_13_mru;
        _zz_cache_tag_3 = ways_3_metas_13_tag;
        _zz_cache_hit_3 = ways_3_metas_13_vld;
        _zz_cache_mru_3 = ways_3_metas_13_mru;
      end
      7'b0001110 : begin
        _zz_cache_tag_0 = ways_0_metas_14_tag;
        _zz_cache_hit_0 = ways_0_metas_14_vld;
        _zz_cache_mru_0 = ways_0_metas_14_mru;
        _zz_cache_tag_1 = ways_1_metas_14_tag;
        _zz_cache_hit_1 = ways_1_metas_14_vld;
        _zz_cache_mru_1 = ways_1_metas_14_mru;
        _zz_cache_tag_2 = ways_2_metas_14_tag;
        _zz_cache_hit_2 = ways_2_metas_14_vld;
        _zz_cache_mru_2 = ways_2_metas_14_mru;
        _zz_cache_tag_3 = ways_3_metas_14_tag;
        _zz_cache_hit_3 = ways_3_metas_14_vld;
        _zz_cache_mru_3 = ways_3_metas_14_mru;
      end
      7'b0001111 : begin
        _zz_cache_tag_0 = ways_0_metas_15_tag;
        _zz_cache_hit_0 = ways_0_metas_15_vld;
        _zz_cache_mru_0 = ways_0_metas_15_mru;
        _zz_cache_tag_1 = ways_1_metas_15_tag;
        _zz_cache_hit_1 = ways_1_metas_15_vld;
        _zz_cache_mru_1 = ways_1_metas_15_mru;
        _zz_cache_tag_2 = ways_2_metas_15_tag;
        _zz_cache_hit_2 = ways_2_metas_15_vld;
        _zz_cache_mru_2 = ways_2_metas_15_mru;
        _zz_cache_tag_3 = ways_3_metas_15_tag;
        _zz_cache_hit_3 = ways_3_metas_15_vld;
        _zz_cache_mru_3 = ways_3_metas_15_mru;
      end
      7'b0010000 : begin
        _zz_cache_tag_0 = ways_0_metas_16_tag;
        _zz_cache_hit_0 = ways_0_metas_16_vld;
        _zz_cache_mru_0 = ways_0_metas_16_mru;
        _zz_cache_tag_1 = ways_1_metas_16_tag;
        _zz_cache_hit_1 = ways_1_metas_16_vld;
        _zz_cache_mru_1 = ways_1_metas_16_mru;
        _zz_cache_tag_2 = ways_2_metas_16_tag;
        _zz_cache_hit_2 = ways_2_metas_16_vld;
        _zz_cache_mru_2 = ways_2_metas_16_mru;
        _zz_cache_tag_3 = ways_3_metas_16_tag;
        _zz_cache_hit_3 = ways_3_metas_16_vld;
        _zz_cache_mru_3 = ways_3_metas_16_mru;
      end
      7'b0010001 : begin
        _zz_cache_tag_0 = ways_0_metas_17_tag;
        _zz_cache_hit_0 = ways_0_metas_17_vld;
        _zz_cache_mru_0 = ways_0_metas_17_mru;
        _zz_cache_tag_1 = ways_1_metas_17_tag;
        _zz_cache_hit_1 = ways_1_metas_17_vld;
        _zz_cache_mru_1 = ways_1_metas_17_mru;
        _zz_cache_tag_2 = ways_2_metas_17_tag;
        _zz_cache_hit_2 = ways_2_metas_17_vld;
        _zz_cache_mru_2 = ways_2_metas_17_mru;
        _zz_cache_tag_3 = ways_3_metas_17_tag;
        _zz_cache_hit_3 = ways_3_metas_17_vld;
        _zz_cache_mru_3 = ways_3_metas_17_mru;
      end
      7'b0010010 : begin
        _zz_cache_tag_0 = ways_0_metas_18_tag;
        _zz_cache_hit_0 = ways_0_metas_18_vld;
        _zz_cache_mru_0 = ways_0_metas_18_mru;
        _zz_cache_tag_1 = ways_1_metas_18_tag;
        _zz_cache_hit_1 = ways_1_metas_18_vld;
        _zz_cache_mru_1 = ways_1_metas_18_mru;
        _zz_cache_tag_2 = ways_2_metas_18_tag;
        _zz_cache_hit_2 = ways_2_metas_18_vld;
        _zz_cache_mru_2 = ways_2_metas_18_mru;
        _zz_cache_tag_3 = ways_3_metas_18_tag;
        _zz_cache_hit_3 = ways_3_metas_18_vld;
        _zz_cache_mru_3 = ways_3_metas_18_mru;
      end
      7'b0010011 : begin
        _zz_cache_tag_0 = ways_0_metas_19_tag;
        _zz_cache_hit_0 = ways_0_metas_19_vld;
        _zz_cache_mru_0 = ways_0_metas_19_mru;
        _zz_cache_tag_1 = ways_1_metas_19_tag;
        _zz_cache_hit_1 = ways_1_metas_19_vld;
        _zz_cache_mru_1 = ways_1_metas_19_mru;
        _zz_cache_tag_2 = ways_2_metas_19_tag;
        _zz_cache_hit_2 = ways_2_metas_19_vld;
        _zz_cache_mru_2 = ways_2_metas_19_mru;
        _zz_cache_tag_3 = ways_3_metas_19_tag;
        _zz_cache_hit_3 = ways_3_metas_19_vld;
        _zz_cache_mru_3 = ways_3_metas_19_mru;
      end
      7'b0010100 : begin
        _zz_cache_tag_0 = ways_0_metas_20_tag;
        _zz_cache_hit_0 = ways_0_metas_20_vld;
        _zz_cache_mru_0 = ways_0_metas_20_mru;
        _zz_cache_tag_1 = ways_1_metas_20_tag;
        _zz_cache_hit_1 = ways_1_metas_20_vld;
        _zz_cache_mru_1 = ways_1_metas_20_mru;
        _zz_cache_tag_2 = ways_2_metas_20_tag;
        _zz_cache_hit_2 = ways_2_metas_20_vld;
        _zz_cache_mru_2 = ways_2_metas_20_mru;
        _zz_cache_tag_3 = ways_3_metas_20_tag;
        _zz_cache_hit_3 = ways_3_metas_20_vld;
        _zz_cache_mru_3 = ways_3_metas_20_mru;
      end
      7'b0010101 : begin
        _zz_cache_tag_0 = ways_0_metas_21_tag;
        _zz_cache_hit_0 = ways_0_metas_21_vld;
        _zz_cache_mru_0 = ways_0_metas_21_mru;
        _zz_cache_tag_1 = ways_1_metas_21_tag;
        _zz_cache_hit_1 = ways_1_metas_21_vld;
        _zz_cache_mru_1 = ways_1_metas_21_mru;
        _zz_cache_tag_2 = ways_2_metas_21_tag;
        _zz_cache_hit_2 = ways_2_metas_21_vld;
        _zz_cache_mru_2 = ways_2_metas_21_mru;
        _zz_cache_tag_3 = ways_3_metas_21_tag;
        _zz_cache_hit_3 = ways_3_metas_21_vld;
        _zz_cache_mru_3 = ways_3_metas_21_mru;
      end
      7'b0010110 : begin
        _zz_cache_tag_0 = ways_0_metas_22_tag;
        _zz_cache_hit_0 = ways_0_metas_22_vld;
        _zz_cache_mru_0 = ways_0_metas_22_mru;
        _zz_cache_tag_1 = ways_1_metas_22_tag;
        _zz_cache_hit_1 = ways_1_metas_22_vld;
        _zz_cache_mru_1 = ways_1_metas_22_mru;
        _zz_cache_tag_2 = ways_2_metas_22_tag;
        _zz_cache_hit_2 = ways_2_metas_22_vld;
        _zz_cache_mru_2 = ways_2_metas_22_mru;
        _zz_cache_tag_3 = ways_3_metas_22_tag;
        _zz_cache_hit_3 = ways_3_metas_22_vld;
        _zz_cache_mru_3 = ways_3_metas_22_mru;
      end
      7'b0010111 : begin
        _zz_cache_tag_0 = ways_0_metas_23_tag;
        _zz_cache_hit_0 = ways_0_metas_23_vld;
        _zz_cache_mru_0 = ways_0_metas_23_mru;
        _zz_cache_tag_1 = ways_1_metas_23_tag;
        _zz_cache_hit_1 = ways_1_metas_23_vld;
        _zz_cache_mru_1 = ways_1_metas_23_mru;
        _zz_cache_tag_2 = ways_2_metas_23_tag;
        _zz_cache_hit_2 = ways_2_metas_23_vld;
        _zz_cache_mru_2 = ways_2_metas_23_mru;
        _zz_cache_tag_3 = ways_3_metas_23_tag;
        _zz_cache_hit_3 = ways_3_metas_23_vld;
        _zz_cache_mru_3 = ways_3_metas_23_mru;
      end
      7'b0011000 : begin
        _zz_cache_tag_0 = ways_0_metas_24_tag;
        _zz_cache_hit_0 = ways_0_metas_24_vld;
        _zz_cache_mru_0 = ways_0_metas_24_mru;
        _zz_cache_tag_1 = ways_1_metas_24_tag;
        _zz_cache_hit_1 = ways_1_metas_24_vld;
        _zz_cache_mru_1 = ways_1_metas_24_mru;
        _zz_cache_tag_2 = ways_2_metas_24_tag;
        _zz_cache_hit_2 = ways_2_metas_24_vld;
        _zz_cache_mru_2 = ways_2_metas_24_mru;
        _zz_cache_tag_3 = ways_3_metas_24_tag;
        _zz_cache_hit_3 = ways_3_metas_24_vld;
        _zz_cache_mru_3 = ways_3_metas_24_mru;
      end
      7'b0011001 : begin
        _zz_cache_tag_0 = ways_0_metas_25_tag;
        _zz_cache_hit_0 = ways_0_metas_25_vld;
        _zz_cache_mru_0 = ways_0_metas_25_mru;
        _zz_cache_tag_1 = ways_1_metas_25_tag;
        _zz_cache_hit_1 = ways_1_metas_25_vld;
        _zz_cache_mru_1 = ways_1_metas_25_mru;
        _zz_cache_tag_2 = ways_2_metas_25_tag;
        _zz_cache_hit_2 = ways_2_metas_25_vld;
        _zz_cache_mru_2 = ways_2_metas_25_mru;
        _zz_cache_tag_3 = ways_3_metas_25_tag;
        _zz_cache_hit_3 = ways_3_metas_25_vld;
        _zz_cache_mru_3 = ways_3_metas_25_mru;
      end
      7'b0011010 : begin
        _zz_cache_tag_0 = ways_0_metas_26_tag;
        _zz_cache_hit_0 = ways_0_metas_26_vld;
        _zz_cache_mru_0 = ways_0_metas_26_mru;
        _zz_cache_tag_1 = ways_1_metas_26_tag;
        _zz_cache_hit_1 = ways_1_metas_26_vld;
        _zz_cache_mru_1 = ways_1_metas_26_mru;
        _zz_cache_tag_2 = ways_2_metas_26_tag;
        _zz_cache_hit_2 = ways_2_metas_26_vld;
        _zz_cache_mru_2 = ways_2_metas_26_mru;
        _zz_cache_tag_3 = ways_3_metas_26_tag;
        _zz_cache_hit_3 = ways_3_metas_26_vld;
        _zz_cache_mru_3 = ways_3_metas_26_mru;
      end
      7'b0011011 : begin
        _zz_cache_tag_0 = ways_0_metas_27_tag;
        _zz_cache_hit_0 = ways_0_metas_27_vld;
        _zz_cache_mru_0 = ways_0_metas_27_mru;
        _zz_cache_tag_1 = ways_1_metas_27_tag;
        _zz_cache_hit_1 = ways_1_metas_27_vld;
        _zz_cache_mru_1 = ways_1_metas_27_mru;
        _zz_cache_tag_2 = ways_2_metas_27_tag;
        _zz_cache_hit_2 = ways_2_metas_27_vld;
        _zz_cache_mru_2 = ways_2_metas_27_mru;
        _zz_cache_tag_3 = ways_3_metas_27_tag;
        _zz_cache_hit_3 = ways_3_metas_27_vld;
        _zz_cache_mru_3 = ways_3_metas_27_mru;
      end
      7'b0011100 : begin
        _zz_cache_tag_0 = ways_0_metas_28_tag;
        _zz_cache_hit_0 = ways_0_metas_28_vld;
        _zz_cache_mru_0 = ways_0_metas_28_mru;
        _zz_cache_tag_1 = ways_1_metas_28_tag;
        _zz_cache_hit_1 = ways_1_metas_28_vld;
        _zz_cache_mru_1 = ways_1_metas_28_mru;
        _zz_cache_tag_2 = ways_2_metas_28_tag;
        _zz_cache_hit_2 = ways_2_metas_28_vld;
        _zz_cache_mru_2 = ways_2_metas_28_mru;
        _zz_cache_tag_3 = ways_3_metas_28_tag;
        _zz_cache_hit_3 = ways_3_metas_28_vld;
        _zz_cache_mru_3 = ways_3_metas_28_mru;
      end
      7'b0011101 : begin
        _zz_cache_tag_0 = ways_0_metas_29_tag;
        _zz_cache_hit_0 = ways_0_metas_29_vld;
        _zz_cache_mru_0 = ways_0_metas_29_mru;
        _zz_cache_tag_1 = ways_1_metas_29_tag;
        _zz_cache_hit_1 = ways_1_metas_29_vld;
        _zz_cache_mru_1 = ways_1_metas_29_mru;
        _zz_cache_tag_2 = ways_2_metas_29_tag;
        _zz_cache_hit_2 = ways_2_metas_29_vld;
        _zz_cache_mru_2 = ways_2_metas_29_mru;
        _zz_cache_tag_3 = ways_3_metas_29_tag;
        _zz_cache_hit_3 = ways_3_metas_29_vld;
        _zz_cache_mru_3 = ways_3_metas_29_mru;
      end
      7'b0011110 : begin
        _zz_cache_tag_0 = ways_0_metas_30_tag;
        _zz_cache_hit_0 = ways_0_metas_30_vld;
        _zz_cache_mru_0 = ways_0_metas_30_mru;
        _zz_cache_tag_1 = ways_1_metas_30_tag;
        _zz_cache_hit_1 = ways_1_metas_30_vld;
        _zz_cache_mru_1 = ways_1_metas_30_mru;
        _zz_cache_tag_2 = ways_2_metas_30_tag;
        _zz_cache_hit_2 = ways_2_metas_30_vld;
        _zz_cache_mru_2 = ways_2_metas_30_mru;
        _zz_cache_tag_3 = ways_3_metas_30_tag;
        _zz_cache_hit_3 = ways_3_metas_30_vld;
        _zz_cache_mru_3 = ways_3_metas_30_mru;
      end
      7'b0011111 : begin
        _zz_cache_tag_0 = ways_0_metas_31_tag;
        _zz_cache_hit_0 = ways_0_metas_31_vld;
        _zz_cache_mru_0 = ways_0_metas_31_mru;
        _zz_cache_tag_1 = ways_1_metas_31_tag;
        _zz_cache_hit_1 = ways_1_metas_31_vld;
        _zz_cache_mru_1 = ways_1_metas_31_mru;
        _zz_cache_tag_2 = ways_2_metas_31_tag;
        _zz_cache_hit_2 = ways_2_metas_31_vld;
        _zz_cache_mru_2 = ways_2_metas_31_mru;
        _zz_cache_tag_3 = ways_3_metas_31_tag;
        _zz_cache_hit_3 = ways_3_metas_31_vld;
        _zz_cache_mru_3 = ways_3_metas_31_mru;
      end
      7'b0100000 : begin
        _zz_cache_tag_0 = ways_0_metas_32_tag;
        _zz_cache_hit_0 = ways_0_metas_32_vld;
        _zz_cache_mru_0 = ways_0_metas_32_mru;
        _zz_cache_tag_1 = ways_1_metas_32_tag;
        _zz_cache_hit_1 = ways_1_metas_32_vld;
        _zz_cache_mru_1 = ways_1_metas_32_mru;
        _zz_cache_tag_2 = ways_2_metas_32_tag;
        _zz_cache_hit_2 = ways_2_metas_32_vld;
        _zz_cache_mru_2 = ways_2_metas_32_mru;
        _zz_cache_tag_3 = ways_3_metas_32_tag;
        _zz_cache_hit_3 = ways_3_metas_32_vld;
        _zz_cache_mru_3 = ways_3_metas_32_mru;
      end
      7'b0100001 : begin
        _zz_cache_tag_0 = ways_0_metas_33_tag;
        _zz_cache_hit_0 = ways_0_metas_33_vld;
        _zz_cache_mru_0 = ways_0_metas_33_mru;
        _zz_cache_tag_1 = ways_1_metas_33_tag;
        _zz_cache_hit_1 = ways_1_metas_33_vld;
        _zz_cache_mru_1 = ways_1_metas_33_mru;
        _zz_cache_tag_2 = ways_2_metas_33_tag;
        _zz_cache_hit_2 = ways_2_metas_33_vld;
        _zz_cache_mru_2 = ways_2_metas_33_mru;
        _zz_cache_tag_3 = ways_3_metas_33_tag;
        _zz_cache_hit_3 = ways_3_metas_33_vld;
        _zz_cache_mru_3 = ways_3_metas_33_mru;
      end
      7'b0100010 : begin
        _zz_cache_tag_0 = ways_0_metas_34_tag;
        _zz_cache_hit_0 = ways_0_metas_34_vld;
        _zz_cache_mru_0 = ways_0_metas_34_mru;
        _zz_cache_tag_1 = ways_1_metas_34_tag;
        _zz_cache_hit_1 = ways_1_metas_34_vld;
        _zz_cache_mru_1 = ways_1_metas_34_mru;
        _zz_cache_tag_2 = ways_2_metas_34_tag;
        _zz_cache_hit_2 = ways_2_metas_34_vld;
        _zz_cache_mru_2 = ways_2_metas_34_mru;
        _zz_cache_tag_3 = ways_3_metas_34_tag;
        _zz_cache_hit_3 = ways_3_metas_34_vld;
        _zz_cache_mru_3 = ways_3_metas_34_mru;
      end
      7'b0100011 : begin
        _zz_cache_tag_0 = ways_0_metas_35_tag;
        _zz_cache_hit_0 = ways_0_metas_35_vld;
        _zz_cache_mru_0 = ways_0_metas_35_mru;
        _zz_cache_tag_1 = ways_1_metas_35_tag;
        _zz_cache_hit_1 = ways_1_metas_35_vld;
        _zz_cache_mru_1 = ways_1_metas_35_mru;
        _zz_cache_tag_2 = ways_2_metas_35_tag;
        _zz_cache_hit_2 = ways_2_metas_35_vld;
        _zz_cache_mru_2 = ways_2_metas_35_mru;
        _zz_cache_tag_3 = ways_3_metas_35_tag;
        _zz_cache_hit_3 = ways_3_metas_35_vld;
        _zz_cache_mru_3 = ways_3_metas_35_mru;
      end
      7'b0100100 : begin
        _zz_cache_tag_0 = ways_0_metas_36_tag;
        _zz_cache_hit_0 = ways_0_metas_36_vld;
        _zz_cache_mru_0 = ways_0_metas_36_mru;
        _zz_cache_tag_1 = ways_1_metas_36_tag;
        _zz_cache_hit_1 = ways_1_metas_36_vld;
        _zz_cache_mru_1 = ways_1_metas_36_mru;
        _zz_cache_tag_2 = ways_2_metas_36_tag;
        _zz_cache_hit_2 = ways_2_metas_36_vld;
        _zz_cache_mru_2 = ways_2_metas_36_mru;
        _zz_cache_tag_3 = ways_3_metas_36_tag;
        _zz_cache_hit_3 = ways_3_metas_36_vld;
        _zz_cache_mru_3 = ways_3_metas_36_mru;
      end
      7'b0100101 : begin
        _zz_cache_tag_0 = ways_0_metas_37_tag;
        _zz_cache_hit_0 = ways_0_metas_37_vld;
        _zz_cache_mru_0 = ways_0_metas_37_mru;
        _zz_cache_tag_1 = ways_1_metas_37_tag;
        _zz_cache_hit_1 = ways_1_metas_37_vld;
        _zz_cache_mru_1 = ways_1_metas_37_mru;
        _zz_cache_tag_2 = ways_2_metas_37_tag;
        _zz_cache_hit_2 = ways_2_metas_37_vld;
        _zz_cache_mru_2 = ways_2_metas_37_mru;
        _zz_cache_tag_3 = ways_3_metas_37_tag;
        _zz_cache_hit_3 = ways_3_metas_37_vld;
        _zz_cache_mru_3 = ways_3_metas_37_mru;
      end
      7'b0100110 : begin
        _zz_cache_tag_0 = ways_0_metas_38_tag;
        _zz_cache_hit_0 = ways_0_metas_38_vld;
        _zz_cache_mru_0 = ways_0_metas_38_mru;
        _zz_cache_tag_1 = ways_1_metas_38_tag;
        _zz_cache_hit_1 = ways_1_metas_38_vld;
        _zz_cache_mru_1 = ways_1_metas_38_mru;
        _zz_cache_tag_2 = ways_2_metas_38_tag;
        _zz_cache_hit_2 = ways_2_metas_38_vld;
        _zz_cache_mru_2 = ways_2_metas_38_mru;
        _zz_cache_tag_3 = ways_3_metas_38_tag;
        _zz_cache_hit_3 = ways_3_metas_38_vld;
        _zz_cache_mru_3 = ways_3_metas_38_mru;
      end
      7'b0100111 : begin
        _zz_cache_tag_0 = ways_0_metas_39_tag;
        _zz_cache_hit_0 = ways_0_metas_39_vld;
        _zz_cache_mru_0 = ways_0_metas_39_mru;
        _zz_cache_tag_1 = ways_1_metas_39_tag;
        _zz_cache_hit_1 = ways_1_metas_39_vld;
        _zz_cache_mru_1 = ways_1_metas_39_mru;
        _zz_cache_tag_2 = ways_2_metas_39_tag;
        _zz_cache_hit_2 = ways_2_metas_39_vld;
        _zz_cache_mru_2 = ways_2_metas_39_mru;
        _zz_cache_tag_3 = ways_3_metas_39_tag;
        _zz_cache_hit_3 = ways_3_metas_39_vld;
        _zz_cache_mru_3 = ways_3_metas_39_mru;
      end
      7'b0101000 : begin
        _zz_cache_tag_0 = ways_0_metas_40_tag;
        _zz_cache_hit_0 = ways_0_metas_40_vld;
        _zz_cache_mru_0 = ways_0_metas_40_mru;
        _zz_cache_tag_1 = ways_1_metas_40_tag;
        _zz_cache_hit_1 = ways_1_metas_40_vld;
        _zz_cache_mru_1 = ways_1_metas_40_mru;
        _zz_cache_tag_2 = ways_2_metas_40_tag;
        _zz_cache_hit_2 = ways_2_metas_40_vld;
        _zz_cache_mru_2 = ways_2_metas_40_mru;
        _zz_cache_tag_3 = ways_3_metas_40_tag;
        _zz_cache_hit_3 = ways_3_metas_40_vld;
        _zz_cache_mru_3 = ways_3_metas_40_mru;
      end
      7'b0101001 : begin
        _zz_cache_tag_0 = ways_0_metas_41_tag;
        _zz_cache_hit_0 = ways_0_metas_41_vld;
        _zz_cache_mru_0 = ways_0_metas_41_mru;
        _zz_cache_tag_1 = ways_1_metas_41_tag;
        _zz_cache_hit_1 = ways_1_metas_41_vld;
        _zz_cache_mru_1 = ways_1_metas_41_mru;
        _zz_cache_tag_2 = ways_2_metas_41_tag;
        _zz_cache_hit_2 = ways_2_metas_41_vld;
        _zz_cache_mru_2 = ways_2_metas_41_mru;
        _zz_cache_tag_3 = ways_3_metas_41_tag;
        _zz_cache_hit_3 = ways_3_metas_41_vld;
        _zz_cache_mru_3 = ways_3_metas_41_mru;
      end
      7'b0101010 : begin
        _zz_cache_tag_0 = ways_0_metas_42_tag;
        _zz_cache_hit_0 = ways_0_metas_42_vld;
        _zz_cache_mru_0 = ways_0_metas_42_mru;
        _zz_cache_tag_1 = ways_1_metas_42_tag;
        _zz_cache_hit_1 = ways_1_metas_42_vld;
        _zz_cache_mru_1 = ways_1_metas_42_mru;
        _zz_cache_tag_2 = ways_2_metas_42_tag;
        _zz_cache_hit_2 = ways_2_metas_42_vld;
        _zz_cache_mru_2 = ways_2_metas_42_mru;
        _zz_cache_tag_3 = ways_3_metas_42_tag;
        _zz_cache_hit_3 = ways_3_metas_42_vld;
        _zz_cache_mru_3 = ways_3_metas_42_mru;
      end
      7'b0101011 : begin
        _zz_cache_tag_0 = ways_0_metas_43_tag;
        _zz_cache_hit_0 = ways_0_metas_43_vld;
        _zz_cache_mru_0 = ways_0_metas_43_mru;
        _zz_cache_tag_1 = ways_1_metas_43_tag;
        _zz_cache_hit_1 = ways_1_metas_43_vld;
        _zz_cache_mru_1 = ways_1_metas_43_mru;
        _zz_cache_tag_2 = ways_2_metas_43_tag;
        _zz_cache_hit_2 = ways_2_metas_43_vld;
        _zz_cache_mru_2 = ways_2_metas_43_mru;
        _zz_cache_tag_3 = ways_3_metas_43_tag;
        _zz_cache_hit_3 = ways_3_metas_43_vld;
        _zz_cache_mru_3 = ways_3_metas_43_mru;
      end
      7'b0101100 : begin
        _zz_cache_tag_0 = ways_0_metas_44_tag;
        _zz_cache_hit_0 = ways_0_metas_44_vld;
        _zz_cache_mru_0 = ways_0_metas_44_mru;
        _zz_cache_tag_1 = ways_1_metas_44_tag;
        _zz_cache_hit_1 = ways_1_metas_44_vld;
        _zz_cache_mru_1 = ways_1_metas_44_mru;
        _zz_cache_tag_2 = ways_2_metas_44_tag;
        _zz_cache_hit_2 = ways_2_metas_44_vld;
        _zz_cache_mru_2 = ways_2_metas_44_mru;
        _zz_cache_tag_3 = ways_3_metas_44_tag;
        _zz_cache_hit_3 = ways_3_metas_44_vld;
        _zz_cache_mru_3 = ways_3_metas_44_mru;
      end
      7'b0101101 : begin
        _zz_cache_tag_0 = ways_0_metas_45_tag;
        _zz_cache_hit_0 = ways_0_metas_45_vld;
        _zz_cache_mru_0 = ways_0_metas_45_mru;
        _zz_cache_tag_1 = ways_1_metas_45_tag;
        _zz_cache_hit_1 = ways_1_metas_45_vld;
        _zz_cache_mru_1 = ways_1_metas_45_mru;
        _zz_cache_tag_2 = ways_2_metas_45_tag;
        _zz_cache_hit_2 = ways_2_metas_45_vld;
        _zz_cache_mru_2 = ways_2_metas_45_mru;
        _zz_cache_tag_3 = ways_3_metas_45_tag;
        _zz_cache_hit_3 = ways_3_metas_45_vld;
        _zz_cache_mru_3 = ways_3_metas_45_mru;
      end
      7'b0101110 : begin
        _zz_cache_tag_0 = ways_0_metas_46_tag;
        _zz_cache_hit_0 = ways_0_metas_46_vld;
        _zz_cache_mru_0 = ways_0_metas_46_mru;
        _zz_cache_tag_1 = ways_1_metas_46_tag;
        _zz_cache_hit_1 = ways_1_metas_46_vld;
        _zz_cache_mru_1 = ways_1_metas_46_mru;
        _zz_cache_tag_2 = ways_2_metas_46_tag;
        _zz_cache_hit_2 = ways_2_metas_46_vld;
        _zz_cache_mru_2 = ways_2_metas_46_mru;
        _zz_cache_tag_3 = ways_3_metas_46_tag;
        _zz_cache_hit_3 = ways_3_metas_46_vld;
        _zz_cache_mru_3 = ways_3_metas_46_mru;
      end
      7'b0101111 : begin
        _zz_cache_tag_0 = ways_0_metas_47_tag;
        _zz_cache_hit_0 = ways_0_metas_47_vld;
        _zz_cache_mru_0 = ways_0_metas_47_mru;
        _zz_cache_tag_1 = ways_1_metas_47_tag;
        _zz_cache_hit_1 = ways_1_metas_47_vld;
        _zz_cache_mru_1 = ways_1_metas_47_mru;
        _zz_cache_tag_2 = ways_2_metas_47_tag;
        _zz_cache_hit_2 = ways_2_metas_47_vld;
        _zz_cache_mru_2 = ways_2_metas_47_mru;
        _zz_cache_tag_3 = ways_3_metas_47_tag;
        _zz_cache_hit_3 = ways_3_metas_47_vld;
        _zz_cache_mru_3 = ways_3_metas_47_mru;
      end
      7'b0110000 : begin
        _zz_cache_tag_0 = ways_0_metas_48_tag;
        _zz_cache_hit_0 = ways_0_metas_48_vld;
        _zz_cache_mru_0 = ways_0_metas_48_mru;
        _zz_cache_tag_1 = ways_1_metas_48_tag;
        _zz_cache_hit_1 = ways_1_metas_48_vld;
        _zz_cache_mru_1 = ways_1_metas_48_mru;
        _zz_cache_tag_2 = ways_2_metas_48_tag;
        _zz_cache_hit_2 = ways_2_metas_48_vld;
        _zz_cache_mru_2 = ways_2_metas_48_mru;
        _zz_cache_tag_3 = ways_3_metas_48_tag;
        _zz_cache_hit_3 = ways_3_metas_48_vld;
        _zz_cache_mru_3 = ways_3_metas_48_mru;
      end
      7'b0110001 : begin
        _zz_cache_tag_0 = ways_0_metas_49_tag;
        _zz_cache_hit_0 = ways_0_metas_49_vld;
        _zz_cache_mru_0 = ways_0_metas_49_mru;
        _zz_cache_tag_1 = ways_1_metas_49_tag;
        _zz_cache_hit_1 = ways_1_metas_49_vld;
        _zz_cache_mru_1 = ways_1_metas_49_mru;
        _zz_cache_tag_2 = ways_2_metas_49_tag;
        _zz_cache_hit_2 = ways_2_metas_49_vld;
        _zz_cache_mru_2 = ways_2_metas_49_mru;
        _zz_cache_tag_3 = ways_3_metas_49_tag;
        _zz_cache_hit_3 = ways_3_metas_49_vld;
        _zz_cache_mru_3 = ways_3_metas_49_mru;
      end
      7'b0110010 : begin
        _zz_cache_tag_0 = ways_0_metas_50_tag;
        _zz_cache_hit_0 = ways_0_metas_50_vld;
        _zz_cache_mru_0 = ways_0_metas_50_mru;
        _zz_cache_tag_1 = ways_1_metas_50_tag;
        _zz_cache_hit_1 = ways_1_metas_50_vld;
        _zz_cache_mru_1 = ways_1_metas_50_mru;
        _zz_cache_tag_2 = ways_2_metas_50_tag;
        _zz_cache_hit_2 = ways_2_metas_50_vld;
        _zz_cache_mru_2 = ways_2_metas_50_mru;
        _zz_cache_tag_3 = ways_3_metas_50_tag;
        _zz_cache_hit_3 = ways_3_metas_50_vld;
        _zz_cache_mru_3 = ways_3_metas_50_mru;
      end
      7'b0110011 : begin
        _zz_cache_tag_0 = ways_0_metas_51_tag;
        _zz_cache_hit_0 = ways_0_metas_51_vld;
        _zz_cache_mru_0 = ways_0_metas_51_mru;
        _zz_cache_tag_1 = ways_1_metas_51_tag;
        _zz_cache_hit_1 = ways_1_metas_51_vld;
        _zz_cache_mru_1 = ways_1_metas_51_mru;
        _zz_cache_tag_2 = ways_2_metas_51_tag;
        _zz_cache_hit_2 = ways_2_metas_51_vld;
        _zz_cache_mru_2 = ways_2_metas_51_mru;
        _zz_cache_tag_3 = ways_3_metas_51_tag;
        _zz_cache_hit_3 = ways_3_metas_51_vld;
        _zz_cache_mru_3 = ways_3_metas_51_mru;
      end
      7'b0110100 : begin
        _zz_cache_tag_0 = ways_0_metas_52_tag;
        _zz_cache_hit_0 = ways_0_metas_52_vld;
        _zz_cache_mru_0 = ways_0_metas_52_mru;
        _zz_cache_tag_1 = ways_1_metas_52_tag;
        _zz_cache_hit_1 = ways_1_metas_52_vld;
        _zz_cache_mru_1 = ways_1_metas_52_mru;
        _zz_cache_tag_2 = ways_2_metas_52_tag;
        _zz_cache_hit_2 = ways_2_metas_52_vld;
        _zz_cache_mru_2 = ways_2_metas_52_mru;
        _zz_cache_tag_3 = ways_3_metas_52_tag;
        _zz_cache_hit_3 = ways_3_metas_52_vld;
        _zz_cache_mru_3 = ways_3_metas_52_mru;
      end
      7'b0110101 : begin
        _zz_cache_tag_0 = ways_0_metas_53_tag;
        _zz_cache_hit_0 = ways_0_metas_53_vld;
        _zz_cache_mru_0 = ways_0_metas_53_mru;
        _zz_cache_tag_1 = ways_1_metas_53_tag;
        _zz_cache_hit_1 = ways_1_metas_53_vld;
        _zz_cache_mru_1 = ways_1_metas_53_mru;
        _zz_cache_tag_2 = ways_2_metas_53_tag;
        _zz_cache_hit_2 = ways_2_metas_53_vld;
        _zz_cache_mru_2 = ways_2_metas_53_mru;
        _zz_cache_tag_3 = ways_3_metas_53_tag;
        _zz_cache_hit_3 = ways_3_metas_53_vld;
        _zz_cache_mru_3 = ways_3_metas_53_mru;
      end
      7'b0110110 : begin
        _zz_cache_tag_0 = ways_0_metas_54_tag;
        _zz_cache_hit_0 = ways_0_metas_54_vld;
        _zz_cache_mru_0 = ways_0_metas_54_mru;
        _zz_cache_tag_1 = ways_1_metas_54_tag;
        _zz_cache_hit_1 = ways_1_metas_54_vld;
        _zz_cache_mru_1 = ways_1_metas_54_mru;
        _zz_cache_tag_2 = ways_2_metas_54_tag;
        _zz_cache_hit_2 = ways_2_metas_54_vld;
        _zz_cache_mru_2 = ways_2_metas_54_mru;
        _zz_cache_tag_3 = ways_3_metas_54_tag;
        _zz_cache_hit_3 = ways_3_metas_54_vld;
        _zz_cache_mru_3 = ways_3_metas_54_mru;
      end
      7'b0110111 : begin
        _zz_cache_tag_0 = ways_0_metas_55_tag;
        _zz_cache_hit_0 = ways_0_metas_55_vld;
        _zz_cache_mru_0 = ways_0_metas_55_mru;
        _zz_cache_tag_1 = ways_1_metas_55_tag;
        _zz_cache_hit_1 = ways_1_metas_55_vld;
        _zz_cache_mru_1 = ways_1_metas_55_mru;
        _zz_cache_tag_2 = ways_2_metas_55_tag;
        _zz_cache_hit_2 = ways_2_metas_55_vld;
        _zz_cache_mru_2 = ways_2_metas_55_mru;
        _zz_cache_tag_3 = ways_3_metas_55_tag;
        _zz_cache_hit_3 = ways_3_metas_55_vld;
        _zz_cache_mru_3 = ways_3_metas_55_mru;
      end
      7'b0111000 : begin
        _zz_cache_tag_0 = ways_0_metas_56_tag;
        _zz_cache_hit_0 = ways_0_metas_56_vld;
        _zz_cache_mru_0 = ways_0_metas_56_mru;
        _zz_cache_tag_1 = ways_1_metas_56_tag;
        _zz_cache_hit_1 = ways_1_metas_56_vld;
        _zz_cache_mru_1 = ways_1_metas_56_mru;
        _zz_cache_tag_2 = ways_2_metas_56_tag;
        _zz_cache_hit_2 = ways_2_metas_56_vld;
        _zz_cache_mru_2 = ways_2_metas_56_mru;
        _zz_cache_tag_3 = ways_3_metas_56_tag;
        _zz_cache_hit_3 = ways_3_metas_56_vld;
        _zz_cache_mru_3 = ways_3_metas_56_mru;
      end
      7'b0111001 : begin
        _zz_cache_tag_0 = ways_0_metas_57_tag;
        _zz_cache_hit_0 = ways_0_metas_57_vld;
        _zz_cache_mru_0 = ways_0_metas_57_mru;
        _zz_cache_tag_1 = ways_1_metas_57_tag;
        _zz_cache_hit_1 = ways_1_metas_57_vld;
        _zz_cache_mru_1 = ways_1_metas_57_mru;
        _zz_cache_tag_2 = ways_2_metas_57_tag;
        _zz_cache_hit_2 = ways_2_metas_57_vld;
        _zz_cache_mru_2 = ways_2_metas_57_mru;
        _zz_cache_tag_3 = ways_3_metas_57_tag;
        _zz_cache_hit_3 = ways_3_metas_57_vld;
        _zz_cache_mru_3 = ways_3_metas_57_mru;
      end
      7'b0111010 : begin
        _zz_cache_tag_0 = ways_0_metas_58_tag;
        _zz_cache_hit_0 = ways_0_metas_58_vld;
        _zz_cache_mru_0 = ways_0_metas_58_mru;
        _zz_cache_tag_1 = ways_1_metas_58_tag;
        _zz_cache_hit_1 = ways_1_metas_58_vld;
        _zz_cache_mru_1 = ways_1_metas_58_mru;
        _zz_cache_tag_2 = ways_2_metas_58_tag;
        _zz_cache_hit_2 = ways_2_metas_58_vld;
        _zz_cache_mru_2 = ways_2_metas_58_mru;
        _zz_cache_tag_3 = ways_3_metas_58_tag;
        _zz_cache_hit_3 = ways_3_metas_58_vld;
        _zz_cache_mru_3 = ways_3_metas_58_mru;
      end
      7'b0111011 : begin
        _zz_cache_tag_0 = ways_0_metas_59_tag;
        _zz_cache_hit_0 = ways_0_metas_59_vld;
        _zz_cache_mru_0 = ways_0_metas_59_mru;
        _zz_cache_tag_1 = ways_1_metas_59_tag;
        _zz_cache_hit_1 = ways_1_metas_59_vld;
        _zz_cache_mru_1 = ways_1_metas_59_mru;
        _zz_cache_tag_2 = ways_2_metas_59_tag;
        _zz_cache_hit_2 = ways_2_metas_59_vld;
        _zz_cache_mru_2 = ways_2_metas_59_mru;
        _zz_cache_tag_3 = ways_3_metas_59_tag;
        _zz_cache_hit_3 = ways_3_metas_59_vld;
        _zz_cache_mru_3 = ways_3_metas_59_mru;
      end
      7'b0111100 : begin
        _zz_cache_tag_0 = ways_0_metas_60_tag;
        _zz_cache_hit_0 = ways_0_metas_60_vld;
        _zz_cache_mru_0 = ways_0_metas_60_mru;
        _zz_cache_tag_1 = ways_1_metas_60_tag;
        _zz_cache_hit_1 = ways_1_metas_60_vld;
        _zz_cache_mru_1 = ways_1_metas_60_mru;
        _zz_cache_tag_2 = ways_2_metas_60_tag;
        _zz_cache_hit_2 = ways_2_metas_60_vld;
        _zz_cache_mru_2 = ways_2_metas_60_mru;
        _zz_cache_tag_3 = ways_3_metas_60_tag;
        _zz_cache_hit_3 = ways_3_metas_60_vld;
        _zz_cache_mru_3 = ways_3_metas_60_mru;
      end
      7'b0111101 : begin
        _zz_cache_tag_0 = ways_0_metas_61_tag;
        _zz_cache_hit_0 = ways_0_metas_61_vld;
        _zz_cache_mru_0 = ways_0_metas_61_mru;
        _zz_cache_tag_1 = ways_1_metas_61_tag;
        _zz_cache_hit_1 = ways_1_metas_61_vld;
        _zz_cache_mru_1 = ways_1_metas_61_mru;
        _zz_cache_tag_2 = ways_2_metas_61_tag;
        _zz_cache_hit_2 = ways_2_metas_61_vld;
        _zz_cache_mru_2 = ways_2_metas_61_mru;
        _zz_cache_tag_3 = ways_3_metas_61_tag;
        _zz_cache_hit_3 = ways_3_metas_61_vld;
        _zz_cache_mru_3 = ways_3_metas_61_mru;
      end
      7'b0111110 : begin
        _zz_cache_tag_0 = ways_0_metas_62_tag;
        _zz_cache_hit_0 = ways_0_metas_62_vld;
        _zz_cache_mru_0 = ways_0_metas_62_mru;
        _zz_cache_tag_1 = ways_1_metas_62_tag;
        _zz_cache_hit_1 = ways_1_metas_62_vld;
        _zz_cache_mru_1 = ways_1_metas_62_mru;
        _zz_cache_tag_2 = ways_2_metas_62_tag;
        _zz_cache_hit_2 = ways_2_metas_62_vld;
        _zz_cache_mru_2 = ways_2_metas_62_mru;
        _zz_cache_tag_3 = ways_3_metas_62_tag;
        _zz_cache_hit_3 = ways_3_metas_62_vld;
        _zz_cache_mru_3 = ways_3_metas_62_mru;
      end
      7'b0111111 : begin
        _zz_cache_tag_0 = ways_0_metas_63_tag;
        _zz_cache_hit_0 = ways_0_metas_63_vld;
        _zz_cache_mru_0 = ways_0_metas_63_mru;
        _zz_cache_tag_1 = ways_1_metas_63_tag;
        _zz_cache_hit_1 = ways_1_metas_63_vld;
        _zz_cache_mru_1 = ways_1_metas_63_mru;
        _zz_cache_tag_2 = ways_2_metas_63_tag;
        _zz_cache_hit_2 = ways_2_metas_63_vld;
        _zz_cache_mru_2 = ways_2_metas_63_mru;
        _zz_cache_tag_3 = ways_3_metas_63_tag;
        _zz_cache_hit_3 = ways_3_metas_63_vld;
        _zz_cache_mru_3 = ways_3_metas_63_mru;
      end
      7'b1000000 : begin
        _zz_cache_tag_0 = ways_0_metas_64_tag;
        _zz_cache_hit_0 = ways_0_metas_64_vld;
        _zz_cache_mru_0 = ways_0_metas_64_mru;
        _zz_cache_tag_1 = ways_1_metas_64_tag;
        _zz_cache_hit_1 = ways_1_metas_64_vld;
        _zz_cache_mru_1 = ways_1_metas_64_mru;
        _zz_cache_tag_2 = ways_2_metas_64_tag;
        _zz_cache_hit_2 = ways_2_metas_64_vld;
        _zz_cache_mru_2 = ways_2_metas_64_mru;
        _zz_cache_tag_3 = ways_3_metas_64_tag;
        _zz_cache_hit_3 = ways_3_metas_64_vld;
        _zz_cache_mru_3 = ways_3_metas_64_mru;
      end
      7'b1000001 : begin
        _zz_cache_tag_0 = ways_0_metas_65_tag;
        _zz_cache_hit_0 = ways_0_metas_65_vld;
        _zz_cache_mru_0 = ways_0_metas_65_mru;
        _zz_cache_tag_1 = ways_1_metas_65_tag;
        _zz_cache_hit_1 = ways_1_metas_65_vld;
        _zz_cache_mru_1 = ways_1_metas_65_mru;
        _zz_cache_tag_2 = ways_2_metas_65_tag;
        _zz_cache_hit_2 = ways_2_metas_65_vld;
        _zz_cache_mru_2 = ways_2_metas_65_mru;
        _zz_cache_tag_3 = ways_3_metas_65_tag;
        _zz_cache_hit_3 = ways_3_metas_65_vld;
        _zz_cache_mru_3 = ways_3_metas_65_mru;
      end
      7'b1000010 : begin
        _zz_cache_tag_0 = ways_0_metas_66_tag;
        _zz_cache_hit_0 = ways_0_metas_66_vld;
        _zz_cache_mru_0 = ways_0_metas_66_mru;
        _zz_cache_tag_1 = ways_1_metas_66_tag;
        _zz_cache_hit_1 = ways_1_metas_66_vld;
        _zz_cache_mru_1 = ways_1_metas_66_mru;
        _zz_cache_tag_2 = ways_2_metas_66_tag;
        _zz_cache_hit_2 = ways_2_metas_66_vld;
        _zz_cache_mru_2 = ways_2_metas_66_mru;
        _zz_cache_tag_3 = ways_3_metas_66_tag;
        _zz_cache_hit_3 = ways_3_metas_66_vld;
        _zz_cache_mru_3 = ways_3_metas_66_mru;
      end
      7'b1000011 : begin
        _zz_cache_tag_0 = ways_0_metas_67_tag;
        _zz_cache_hit_0 = ways_0_metas_67_vld;
        _zz_cache_mru_0 = ways_0_metas_67_mru;
        _zz_cache_tag_1 = ways_1_metas_67_tag;
        _zz_cache_hit_1 = ways_1_metas_67_vld;
        _zz_cache_mru_1 = ways_1_metas_67_mru;
        _zz_cache_tag_2 = ways_2_metas_67_tag;
        _zz_cache_hit_2 = ways_2_metas_67_vld;
        _zz_cache_mru_2 = ways_2_metas_67_mru;
        _zz_cache_tag_3 = ways_3_metas_67_tag;
        _zz_cache_hit_3 = ways_3_metas_67_vld;
        _zz_cache_mru_3 = ways_3_metas_67_mru;
      end
      7'b1000100 : begin
        _zz_cache_tag_0 = ways_0_metas_68_tag;
        _zz_cache_hit_0 = ways_0_metas_68_vld;
        _zz_cache_mru_0 = ways_0_metas_68_mru;
        _zz_cache_tag_1 = ways_1_metas_68_tag;
        _zz_cache_hit_1 = ways_1_metas_68_vld;
        _zz_cache_mru_1 = ways_1_metas_68_mru;
        _zz_cache_tag_2 = ways_2_metas_68_tag;
        _zz_cache_hit_2 = ways_2_metas_68_vld;
        _zz_cache_mru_2 = ways_2_metas_68_mru;
        _zz_cache_tag_3 = ways_3_metas_68_tag;
        _zz_cache_hit_3 = ways_3_metas_68_vld;
        _zz_cache_mru_3 = ways_3_metas_68_mru;
      end
      7'b1000101 : begin
        _zz_cache_tag_0 = ways_0_metas_69_tag;
        _zz_cache_hit_0 = ways_0_metas_69_vld;
        _zz_cache_mru_0 = ways_0_metas_69_mru;
        _zz_cache_tag_1 = ways_1_metas_69_tag;
        _zz_cache_hit_1 = ways_1_metas_69_vld;
        _zz_cache_mru_1 = ways_1_metas_69_mru;
        _zz_cache_tag_2 = ways_2_metas_69_tag;
        _zz_cache_hit_2 = ways_2_metas_69_vld;
        _zz_cache_mru_2 = ways_2_metas_69_mru;
        _zz_cache_tag_3 = ways_3_metas_69_tag;
        _zz_cache_hit_3 = ways_3_metas_69_vld;
        _zz_cache_mru_3 = ways_3_metas_69_mru;
      end
      7'b1000110 : begin
        _zz_cache_tag_0 = ways_0_metas_70_tag;
        _zz_cache_hit_0 = ways_0_metas_70_vld;
        _zz_cache_mru_0 = ways_0_metas_70_mru;
        _zz_cache_tag_1 = ways_1_metas_70_tag;
        _zz_cache_hit_1 = ways_1_metas_70_vld;
        _zz_cache_mru_1 = ways_1_metas_70_mru;
        _zz_cache_tag_2 = ways_2_metas_70_tag;
        _zz_cache_hit_2 = ways_2_metas_70_vld;
        _zz_cache_mru_2 = ways_2_metas_70_mru;
        _zz_cache_tag_3 = ways_3_metas_70_tag;
        _zz_cache_hit_3 = ways_3_metas_70_vld;
        _zz_cache_mru_3 = ways_3_metas_70_mru;
      end
      7'b1000111 : begin
        _zz_cache_tag_0 = ways_0_metas_71_tag;
        _zz_cache_hit_0 = ways_0_metas_71_vld;
        _zz_cache_mru_0 = ways_0_metas_71_mru;
        _zz_cache_tag_1 = ways_1_metas_71_tag;
        _zz_cache_hit_1 = ways_1_metas_71_vld;
        _zz_cache_mru_1 = ways_1_metas_71_mru;
        _zz_cache_tag_2 = ways_2_metas_71_tag;
        _zz_cache_hit_2 = ways_2_metas_71_vld;
        _zz_cache_mru_2 = ways_2_metas_71_mru;
        _zz_cache_tag_3 = ways_3_metas_71_tag;
        _zz_cache_hit_3 = ways_3_metas_71_vld;
        _zz_cache_mru_3 = ways_3_metas_71_mru;
      end
      7'b1001000 : begin
        _zz_cache_tag_0 = ways_0_metas_72_tag;
        _zz_cache_hit_0 = ways_0_metas_72_vld;
        _zz_cache_mru_0 = ways_0_metas_72_mru;
        _zz_cache_tag_1 = ways_1_metas_72_tag;
        _zz_cache_hit_1 = ways_1_metas_72_vld;
        _zz_cache_mru_1 = ways_1_metas_72_mru;
        _zz_cache_tag_2 = ways_2_metas_72_tag;
        _zz_cache_hit_2 = ways_2_metas_72_vld;
        _zz_cache_mru_2 = ways_2_metas_72_mru;
        _zz_cache_tag_3 = ways_3_metas_72_tag;
        _zz_cache_hit_3 = ways_3_metas_72_vld;
        _zz_cache_mru_3 = ways_3_metas_72_mru;
      end
      7'b1001001 : begin
        _zz_cache_tag_0 = ways_0_metas_73_tag;
        _zz_cache_hit_0 = ways_0_metas_73_vld;
        _zz_cache_mru_0 = ways_0_metas_73_mru;
        _zz_cache_tag_1 = ways_1_metas_73_tag;
        _zz_cache_hit_1 = ways_1_metas_73_vld;
        _zz_cache_mru_1 = ways_1_metas_73_mru;
        _zz_cache_tag_2 = ways_2_metas_73_tag;
        _zz_cache_hit_2 = ways_2_metas_73_vld;
        _zz_cache_mru_2 = ways_2_metas_73_mru;
        _zz_cache_tag_3 = ways_3_metas_73_tag;
        _zz_cache_hit_3 = ways_3_metas_73_vld;
        _zz_cache_mru_3 = ways_3_metas_73_mru;
      end
      7'b1001010 : begin
        _zz_cache_tag_0 = ways_0_metas_74_tag;
        _zz_cache_hit_0 = ways_0_metas_74_vld;
        _zz_cache_mru_0 = ways_0_metas_74_mru;
        _zz_cache_tag_1 = ways_1_metas_74_tag;
        _zz_cache_hit_1 = ways_1_metas_74_vld;
        _zz_cache_mru_1 = ways_1_metas_74_mru;
        _zz_cache_tag_2 = ways_2_metas_74_tag;
        _zz_cache_hit_2 = ways_2_metas_74_vld;
        _zz_cache_mru_2 = ways_2_metas_74_mru;
        _zz_cache_tag_3 = ways_3_metas_74_tag;
        _zz_cache_hit_3 = ways_3_metas_74_vld;
        _zz_cache_mru_3 = ways_3_metas_74_mru;
      end
      7'b1001011 : begin
        _zz_cache_tag_0 = ways_0_metas_75_tag;
        _zz_cache_hit_0 = ways_0_metas_75_vld;
        _zz_cache_mru_0 = ways_0_metas_75_mru;
        _zz_cache_tag_1 = ways_1_metas_75_tag;
        _zz_cache_hit_1 = ways_1_metas_75_vld;
        _zz_cache_mru_1 = ways_1_metas_75_mru;
        _zz_cache_tag_2 = ways_2_metas_75_tag;
        _zz_cache_hit_2 = ways_2_metas_75_vld;
        _zz_cache_mru_2 = ways_2_metas_75_mru;
        _zz_cache_tag_3 = ways_3_metas_75_tag;
        _zz_cache_hit_3 = ways_3_metas_75_vld;
        _zz_cache_mru_3 = ways_3_metas_75_mru;
      end
      7'b1001100 : begin
        _zz_cache_tag_0 = ways_0_metas_76_tag;
        _zz_cache_hit_0 = ways_0_metas_76_vld;
        _zz_cache_mru_0 = ways_0_metas_76_mru;
        _zz_cache_tag_1 = ways_1_metas_76_tag;
        _zz_cache_hit_1 = ways_1_metas_76_vld;
        _zz_cache_mru_1 = ways_1_metas_76_mru;
        _zz_cache_tag_2 = ways_2_metas_76_tag;
        _zz_cache_hit_2 = ways_2_metas_76_vld;
        _zz_cache_mru_2 = ways_2_metas_76_mru;
        _zz_cache_tag_3 = ways_3_metas_76_tag;
        _zz_cache_hit_3 = ways_3_metas_76_vld;
        _zz_cache_mru_3 = ways_3_metas_76_mru;
      end
      7'b1001101 : begin
        _zz_cache_tag_0 = ways_0_metas_77_tag;
        _zz_cache_hit_0 = ways_0_metas_77_vld;
        _zz_cache_mru_0 = ways_0_metas_77_mru;
        _zz_cache_tag_1 = ways_1_metas_77_tag;
        _zz_cache_hit_1 = ways_1_metas_77_vld;
        _zz_cache_mru_1 = ways_1_metas_77_mru;
        _zz_cache_tag_2 = ways_2_metas_77_tag;
        _zz_cache_hit_2 = ways_2_metas_77_vld;
        _zz_cache_mru_2 = ways_2_metas_77_mru;
        _zz_cache_tag_3 = ways_3_metas_77_tag;
        _zz_cache_hit_3 = ways_3_metas_77_vld;
        _zz_cache_mru_3 = ways_3_metas_77_mru;
      end
      7'b1001110 : begin
        _zz_cache_tag_0 = ways_0_metas_78_tag;
        _zz_cache_hit_0 = ways_0_metas_78_vld;
        _zz_cache_mru_0 = ways_0_metas_78_mru;
        _zz_cache_tag_1 = ways_1_metas_78_tag;
        _zz_cache_hit_1 = ways_1_metas_78_vld;
        _zz_cache_mru_1 = ways_1_metas_78_mru;
        _zz_cache_tag_2 = ways_2_metas_78_tag;
        _zz_cache_hit_2 = ways_2_metas_78_vld;
        _zz_cache_mru_2 = ways_2_metas_78_mru;
        _zz_cache_tag_3 = ways_3_metas_78_tag;
        _zz_cache_hit_3 = ways_3_metas_78_vld;
        _zz_cache_mru_3 = ways_3_metas_78_mru;
      end
      7'b1001111 : begin
        _zz_cache_tag_0 = ways_0_metas_79_tag;
        _zz_cache_hit_0 = ways_0_metas_79_vld;
        _zz_cache_mru_0 = ways_0_metas_79_mru;
        _zz_cache_tag_1 = ways_1_metas_79_tag;
        _zz_cache_hit_1 = ways_1_metas_79_vld;
        _zz_cache_mru_1 = ways_1_metas_79_mru;
        _zz_cache_tag_2 = ways_2_metas_79_tag;
        _zz_cache_hit_2 = ways_2_metas_79_vld;
        _zz_cache_mru_2 = ways_2_metas_79_mru;
        _zz_cache_tag_3 = ways_3_metas_79_tag;
        _zz_cache_hit_3 = ways_3_metas_79_vld;
        _zz_cache_mru_3 = ways_3_metas_79_mru;
      end
      7'b1010000 : begin
        _zz_cache_tag_0 = ways_0_metas_80_tag;
        _zz_cache_hit_0 = ways_0_metas_80_vld;
        _zz_cache_mru_0 = ways_0_metas_80_mru;
        _zz_cache_tag_1 = ways_1_metas_80_tag;
        _zz_cache_hit_1 = ways_1_metas_80_vld;
        _zz_cache_mru_1 = ways_1_metas_80_mru;
        _zz_cache_tag_2 = ways_2_metas_80_tag;
        _zz_cache_hit_2 = ways_2_metas_80_vld;
        _zz_cache_mru_2 = ways_2_metas_80_mru;
        _zz_cache_tag_3 = ways_3_metas_80_tag;
        _zz_cache_hit_3 = ways_3_metas_80_vld;
        _zz_cache_mru_3 = ways_3_metas_80_mru;
      end
      7'b1010001 : begin
        _zz_cache_tag_0 = ways_0_metas_81_tag;
        _zz_cache_hit_0 = ways_0_metas_81_vld;
        _zz_cache_mru_0 = ways_0_metas_81_mru;
        _zz_cache_tag_1 = ways_1_metas_81_tag;
        _zz_cache_hit_1 = ways_1_metas_81_vld;
        _zz_cache_mru_1 = ways_1_metas_81_mru;
        _zz_cache_tag_2 = ways_2_metas_81_tag;
        _zz_cache_hit_2 = ways_2_metas_81_vld;
        _zz_cache_mru_2 = ways_2_metas_81_mru;
        _zz_cache_tag_3 = ways_3_metas_81_tag;
        _zz_cache_hit_3 = ways_3_metas_81_vld;
        _zz_cache_mru_3 = ways_3_metas_81_mru;
      end
      7'b1010010 : begin
        _zz_cache_tag_0 = ways_0_metas_82_tag;
        _zz_cache_hit_0 = ways_0_metas_82_vld;
        _zz_cache_mru_0 = ways_0_metas_82_mru;
        _zz_cache_tag_1 = ways_1_metas_82_tag;
        _zz_cache_hit_1 = ways_1_metas_82_vld;
        _zz_cache_mru_1 = ways_1_metas_82_mru;
        _zz_cache_tag_2 = ways_2_metas_82_tag;
        _zz_cache_hit_2 = ways_2_metas_82_vld;
        _zz_cache_mru_2 = ways_2_metas_82_mru;
        _zz_cache_tag_3 = ways_3_metas_82_tag;
        _zz_cache_hit_3 = ways_3_metas_82_vld;
        _zz_cache_mru_3 = ways_3_metas_82_mru;
      end
      7'b1010011 : begin
        _zz_cache_tag_0 = ways_0_metas_83_tag;
        _zz_cache_hit_0 = ways_0_metas_83_vld;
        _zz_cache_mru_0 = ways_0_metas_83_mru;
        _zz_cache_tag_1 = ways_1_metas_83_tag;
        _zz_cache_hit_1 = ways_1_metas_83_vld;
        _zz_cache_mru_1 = ways_1_metas_83_mru;
        _zz_cache_tag_2 = ways_2_metas_83_tag;
        _zz_cache_hit_2 = ways_2_metas_83_vld;
        _zz_cache_mru_2 = ways_2_metas_83_mru;
        _zz_cache_tag_3 = ways_3_metas_83_tag;
        _zz_cache_hit_3 = ways_3_metas_83_vld;
        _zz_cache_mru_3 = ways_3_metas_83_mru;
      end
      7'b1010100 : begin
        _zz_cache_tag_0 = ways_0_metas_84_tag;
        _zz_cache_hit_0 = ways_0_metas_84_vld;
        _zz_cache_mru_0 = ways_0_metas_84_mru;
        _zz_cache_tag_1 = ways_1_metas_84_tag;
        _zz_cache_hit_1 = ways_1_metas_84_vld;
        _zz_cache_mru_1 = ways_1_metas_84_mru;
        _zz_cache_tag_2 = ways_2_metas_84_tag;
        _zz_cache_hit_2 = ways_2_metas_84_vld;
        _zz_cache_mru_2 = ways_2_metas_84_mru;
        _zz_cache_tag_3 = ways_3_metas_84_tag;
        _zz_cache_hit_3 = ways_3_metas_84_vld;
        _zz_cache_mru_3 = ways_3_metas_84_mru;
      end
      7'b1010101 : begin
        _zz_cache_tag_0 = ways_0_metas_85_tag;
        _zz_cache_hit_0 = ways_0_metas_85_vld;
        _zz_cache_mru_0 = ways_0_metas_85_mru;
        _zz_cache_tag_1 = ways_1_metas_85_tag;
        _zz_cache_hit_1 = ways_1_metas_85_vld;
        _zz_cache_mru_1 = ways_1_metas_85_mru;
        _zz_cache_tag_2 = ways_2_metas_85_tag;
        _zz_cache_hit_2 = ways_2_metas_85_vld;
        _zz_cache_mru_2 = ways_2_metas_85_mru;
        _zz_cache_tag_3 = ways_3_metas_85_tag;
        _zz_cache_hit_3 = ways_3_metas_85_vld;
        _zz_cache_mru_3 = ways_3_metas_85_mru;
      end
      7'b1010110 : begin
        _zz_cache_tag_0 = ways_0_metas_86_tag;
        _zz_cache_hit_0 = ways_0_metas_86_vld;
        _zz_cache_mru_0 = ways_0_metas_86_mru;
        _zz_cache_tag_1 = ways_1_metas_86_tag;
        _zz_cache_hit_1 = ways_1_metas_86_vld;
        _zz_cache_mru_1 = ways_1_metas_86_mru;
        _zz_cache_tag_2 = ways_2_metas_86_tag;
        _zz_cache_hit_2 = ways_2_metas_86_vld;
        _zz_cache_mru_2 = ways_2_metas_86_mru;
        _zz_cache_tag_3 = ways_3_metas_86_tag;
        _zz_cache_hit_3 = ways_3_metas_86_vld;
        _zz_cache_mru_3 = ways_3_metas_86_mru;
      end
      7'b1010111 : begin
        _zz_cache_tag_0 = ways_0_metas_87_tag;
        _zz_cache_hit_0 = ways_0_metas_87_vld;
        _zz_cache_mru_0 = ways_0_metas_87_mru;
        _zz_cache_tag_1 = ways_1_metas_87_tag;
        _zz_cache_hit_1 = ways_1_metas_87_vld;
        _zz_cache_mru_1 = ways_1_metas_87_mru;
        _zz_cache_tag_2 = ways_2_metas_87_tag;
        _zz_cache_hit_2 = ways_2_metas_87_vld;
        _zz_cache_mru_2 = ways_2_metas_87_mru;
        _zz_cache_tag_3 = ways_3_metas_87_tag;
        _zz_cache_hit_3 = ways_3_metas_87_vld;
        _zz_cache_mru_3 = ways_3_metas_87_mru;
      end
      7'b1011000 : begin
        _zz_cache_tag_0 = ways_0_metas_88_tag;
        _zz_cache_hit_0 = ways_0_metas_88_vld;
        _zz_cache_mru_0 = ways_0_metas_88_mru;
        _zz_cache_tag_1 = ways_1_metas_88_tag;
        _zz_cache_hit_1 = ways_1_metas_88_vld;
        _zz_cache_mru_1 = ways_1_metas_88_mru;
        _zz_cache_tag_2 = ways_2_metas_88_tag;
        _zz_cache_hit_2 = ways_2_metas_88_vld;
        _zz_cache_mru_2 = ways_2_metas_88_mru;
        _zz_cache_tag_3 = ways_3_metas_88_tag;
        _zz_cache_hit_3 = ways_3_metas_88_vld;
        _zz_cache_mru_3 = ways_3_metas_88_mru;
      end
      7'b1011001 : begin
        _zz_cache_tag_0 = ways_0_metas_89_tag;
        _zz_cache_hit_0 = ways_0_metas_89_vld;
        _zz_cache_mru_0 = ways_0_metas_89_mru;
        _zz_cache_tag_1 = ways_1_metas_89_tag;
        _zz_cache_hit_1 = ways_1_metas_89_vld;
        _zz_cache_mru_1 = ways_1_metas_89_mru;
        _zz_cache_tag_2 = ways_2_metas_89_tag;
        _zz_cache_hit_2 = ways_2_metas_89_vld;
        _zz_cache_mru_2 = ways_2_metas_89_mru;
        _zz_cache_tag_3 = ways_3_metas_89_tag;
        _zz_cache_hit_3 = ways_3_metas_89_vld;
        _zz_cache_mru_3 = ways_3_metas_89_mru;
      end
      7'b1011010 : begin
        _zz_cache_tag_0 = ways_0_metas_90_tag;
        _zz_cache_hit_0 = ways_0_metas_90_vld;
        _zz_cache_mru_0 = ways_0_metas_90_mru;
        _zz_cache_tag_1 = ways_1_metas_90_tag;
        _zz_cache_hit_1 = ways_1_metas_90_vld;
        _zz_cache_mru_1 = ways_1_metas_90_mru;
        _zz_cache_tag_2 = ways_2_metas_90_tag;
        _zz_cache_hit_2 = ways_2_metas_90_vld;
        _zz_cache_mru_2 = ways_2_metas_90_mru;
        _zz_cache_tag_3 = ways_3_metas_90_tag;
        _zz_cache_hit_3 = ways_3_metas_90_vld;
        _zz_cache_mru_3 = ways_3_metas_90_mru;
      end
      7'b1011011 : begin
        _zz_cache_tag_0 = ways_0_metas_91_tag;
        _zz_cache_hit_0 = ways_0_metas_91_vld;
        _zz_cache_mru_0 = ways_0_metas_91_mru;
        _zz_cache_tag_1 = ways_1_metas_91_tag;
        _zz_cache_hit_1 = ways_1_metas_91_vld;
        _zz_cache_mru_1 = ways_1_metas_91_mru;
        _zz_cache_tag_2 = ways_2_metas_91_tag;
        _zz_cache_hit_2 = ways_2_metas_91_vld;
        _zz_cache_mru_2 = ways_2_metas_91_mru;
        _zz_cache_tag_3 = ways_3_metas_91_tag;
        _zz_cache_hit_3 = ways_3_metas_91_vld;
        _zz_cache_mru_3 = ways_3_metas_91_mru;
      end
      7'b1011100 : begin
        _zz_cache_tag_0 = ways_0_metas_92_tag;
        _zz_cache_hit_0 = ways_0_metas_92_vld;
        _zz_cache_mru_0 = ways_0_metas_92_mru;
        _zz_cache_tag_1 = ways_1_metas_92_tag;
        _zz_cache_hit_1 = ways_1_metas_92_vld;
        _zz_cache_mru_1 = ways_1_metas_92_mru;
        _zz_cache_tag_2 = ways_2_metas_92_tag;
        _zz_cache_hit_2 = ways_2_metas_92_vld;
        _zz_cache_mru_2 = ways_2_metas_92_mru;
        _zz_cache_tag_3 = ways_3_metas_92_tag;
        _zz_cache_hit_3 = ways_3_metas_92_vld;
        _zz_cache_mru_3 = ways_3_metas_92_mru;
      end
      7'b1011101 : begin
        _zz_cache_tag_0 = ways_0_metas_93_tag;
        _zz_cache_hit_0 = ways_0_metas_93_vld;
        _zz_cache_mru_0 = ways_0_metas_93_mru;
        _zz_cache_tag_1 = ways_1_metas_93_tag;
        _zz_cache_hit_1 = ways_1_metas_93_vld;
        _zz_cache_mru_1 = ways_1_metas_93_mru;
        _zz_cache_tag_2 = ways_2_metas_93_tag;
        _zz_cache_hit_2 = ways_2_metas_93_vld;
        _zz_cache_mru_2 = ways_2_metas_93_mru;
        _zz_cache_tag_3 = ways_3_metas_93_tag;
        _zz_cache_hit_3 = ways_3_metas_93_vld;
        _zz_cache_mru_3 = ways_3_metas_93_mru;
      end
      7'b1011110 : begin
        _zz_cache_tag_0 = ways_0_metas_94_tag;
        _zz_cache_hit_0 = ways_0_metas_94_vld;
        _zz_cache_mru_0 = ways_0_metas_94_mru;
        _zz_cache_tag_1 = ways_1_metas_94_tag;
        _zz_cache_hit_1 = ways_1_metas_94_vld;
        _zz_cache_mru_1 = ways_1_metas_94_mru;
        _zz_cache_tag_2 = ways_2_metas_94_tag;
        _zz_cache_hit_2 = ways_2_metas_94_vld;
        _zz_cache_mru_2 = ways_2_metas_94_mru;
        _zz_cache_tag_3 = ways_3_metas_94_tag;
        _zz_cache_hit_3 = ways_3_metas_94_vld;
        _zz_cache_mru_3 = ways_3_metas_94_mru;
      end
      7'b1011111 : begin
        _zz_cache_tag_0 = ways_0_metas_95_tag;
        _zz_cache_hit_0 = ways_0_metas_95_vld;
        _zz_cache_mru_0 = ways_0_metas_95_mru;
        _zz_cache_tag_1 = ways_1_metas_95_tag;
        _zz_cache_hit_1 = ways_1_metas_95_vld;
        _zz_cache_mru_1 = ways_1_metas_95_mru;
        _zz_cache_tag_2 = ways_2_metas_95_tag;
        _zz_cache_hit_2 = ways_2_metas_95_vld;
        _zz_cache_mru_2 = ways_2_metas_95_mru;
        _zz_cache_tag_3 = ways_3_metas_95_tag;
        _zz_cache_hit_3 = ways_3_metas_95_vld;
        _zz_cache_mru_3 = ways_3_metas_95_mru;
      end
      7'b1100000 : begin
        _zz_cache_tag_0 = ways_0_metas_96_tag;
        _zz_cache_hit_0 = ways_0_metas_96_vld;
        _zz_cache_mru_0 = ways_0_metas_96_mru;
        _zz_cache_tag_1 = ways_1_metas_96_tag;
        _zz_cache_hit_1 = ways_1_metas_96_vld;
        _zz_cache_mru_1 = ways_1_metas_96_mru;
        _zz_cache_tag_2 = ways_2_metas_96_tag;
        _zz_cache_hit_2 = ways_2_metas_96_vld;
        _zz_cache_mru_2 = ways_2_metas_96_mru;
        _zz_cache_tag_3 = ways_3_metas_96_tag;
        _zz_cache_hit_3 = ways_3_metas_96_vld;
        _zz_cache_mru_3 = ways_3_metas_96_mru;
      end
      7'b1100001 : begin
        _zz_cache_tag_0 = ways_0_metas_97_tag;
        _zz_cache_hit_0 = ways_0_metas_97_vld;
        _zz_cache_mru_0 = ways_0_metas_97_mru;
        _zz_cache_tag_1 = ways_1_metas_97_tag;
        _zz_cache_hit_1 = ways_1_metas_97_vld;
        _zz_cache_mru_1 = ways_1_metas_97_mru;
        _zz_cache_tag_2 = ways_2_metas_97_tag;
        _zz_cache_hit_2 = ways_2_metas_97_vld;
        _zz_cache_mru_2 = ways_2_metas_97_mru;
        _zz_cache_tag_3 = ways_3_metas_97_tag;
        _zz_cache_hit_3 = ways_3_metas_97_vld;
        _zz_cache_mru_3 = ways_3_metas_97_mru;
      end
      7'b1100010 : begin
        _zz_cache_tag_0 = ways_0_metas_98_tag;
        _zz_cache_hit_0 = ways_0_metas_98_vld;
        _zz_cache_mru_0 = ways_0_metas_98_mru;
        _zz_cache_tag_1 = ways_1_metas_98_tag;
        _zz_cache_hit_1 = ways_1_metas_98_vld;
        _zz_cache_mru_1 = ways_1_metas_98_mru;
        _zz_cache_tag_2 = ways_2_metas_98_tag;
        _zz_cache_hit_2 = ways_2_metas_98_vld;
        _zz_cache_mru_2 = ways_2_metas_98_mru;
        _zz_cache_tag_3 = ways_3_metas_98_tag;
        _zz_cache_hit_3 = ways_3_metas_98_vld;
        _zz_cache_mru_3 = ways_3_metas_98_mru;
      end
      7'b1100011 : begin
        _zz_cache_tag_0 = ways_0_metas_99_tag;
        _zz_cache_hit_0 = ways_0_metas_99_vld;
        _zz_cache_mru_0 = ways_0_metas_99_mru;
        _zz_cache_tag_1 = ways_1_metas_99_tag;
        _zz_cache_hit_1 = ways_1_metas_99_vld;
        _zz_cache_mru_1 = ways_1_metas_99_mru;
        _zz_cache_tag_2 = ways_2_metas_99_tag;
        _zz_cache_hit_2 = ways_2_metas_99_vld;
        _zz_cache_mru_2 = ways_2_metas_99_mru;
        _zz_cache_tag_3 = ways_3_metas_99_tag;
        _zz_cache_hit_3 = ways_3_metas_99_vld;
        _zz_cache_mru_3 = ways_3_metas_99_mru;
      end
      7'b1100100 : begin
        _zz_cache_tag_0 = ways_0_metas_100_tag;
        _zz_cache_hit_0 = ways_0_metas_100_vld;
        _zz_cache_mru_0 = ways_0_metas_100_mru;
        _zz_cache_tag_1 = ways_1_metas_100_tag;
        _zz_cache_hit_1 = ways_1_metas_100_vld;
        _zz_cache_mru_1 = ways_1_metas_100_mru;
        _zz_cache_tag_2 = ways_2_metas_100_tag;
        _zz_cache_hit_2 = ways_2_metas_100_vld;
        _zz_cache_mru_2 = ways_2_metas_100_mru;
        _zz_cache_tag_3 = ways_3_metas_100_tag;
        _zz_cache_hit_3 = ways_3_metas_100_vld;
        _zz_cache_mru_3 = ways_3_metas_100_mru;
      end
      7'b1100101 : begin
        _zz_cache_tag_0 = ways_0_metas_101_tag;
        _zz_cache_hit_0 = ways_0_metas_101_vld;
        _zz_cache_mru_0 = ways_0_metas_101_mru;
        _zz_cache_tag_1 = ways_1_metas_101_tag;
        _zz_cache_hit_1 = ways_1_metas_101_vld;
        _zz_cache_mru_1 = ways_1_metas_101_mru;
        _zz_cache_tag_2 = ways_2_metas_101_tag;
        _zz_cache_hit_2 = ways_2_metas_101_vld;
        _zz_cache_mru_2 = ways_2_metas_101_mru;
        _zz_cache_tag_3 = ways_3_metas_101_tag;
        _zz_cache_hit_3 = ways_3_metas_101_vld;
        _zz_cache_mru_3 = ways_3_metas_101_mru;
      end
      7'b1100110 : begin
        _zz_cache_tag_0 = ways_0_metas_102_tag;
        _zz_cache_hit_0 = ways_0_metas_102_vld;
        _zz_cache_mru_0 = ways_0_metas_102_mru;
        _zz_cache_tag_1 = ways_1_metas_102_tag;
        _zz_cache_hit_1 = ways_1_metas_102_vld;
        _zz_cache_mru_1 = ways_1_metas_102_mru;
        _zz_cache_tag_2 = ways_2_metas_102_tag;
        _zz_cache_hit_2 = ways_2_metas_102_vld;
        _zz_cache_mru_2 = ways_2_metas_102_mru;
        _zz_cache_tag_3 = ways_3_metas_102_tag;
        _zz_cache_hit_3 = ways_3_metas_102_vld;
        _zz_cache_mru_3 = ways_3_metas_102_mru;
      end
      7'b1100111 : begin
        _zz_cache_tag_0 = ways_0_metas_103_tag;
        _zz_cache_hit_0 = ways_0_metas_103_vld;
        _zz_cache_mru_0 = ways_0_metas_103_mru;
        _zz_cache_tag_1 = ways_1_metas_103_tag;
        _zz_cache_hit_1 = ways_1_metas_103_vld;
        _zz_cache_mru_1 = ways_1_metas_103_mru;
        _zz_cache_tag_2 = ways_2_metas_103_tag;
        _zz_cache_hit_2 = ways_2_metas_103_vld;
        _zz_cache_mru_2 = ways_2_metas_103_mru;
        _zz_cache_tag_3 = ways_3_metas_103_tag;
        _zz_cache_hit_3 = ways_3_metas_103_vld;
        _zz_cache_mru_3 = ways_3_metas_103_mru;
      end
      7'b1101000 : begin
        _zz_cache_tag_0 = ways_0_metas_104_tag;
        _zz_cache_hit_0 = ways_0_metas_104_vld;
        _zz_cache_mru_0 = ways_0_metas_104_mru;
        _zz_cache_tag_1 = ways_1_metas_104_tag;
        _zz_cache_hit_1 = ways_1_metas_104_vld;
        _zz_cache_mru_1 = ways_1_metas_104_mru;
        _zz_cache_tag_2 = ways_2_metas_104_tag;
        _zz_cache_hit_2 = ways_2_metas_104_vld;
        _zz_cache_mru_2 = ways_2_metas_104_mru;
        _zz_cache_tag_3 = ways_3_metas_104_tag;
        _zz_cache_hit_3 = ways_3_metas_104_vld;
        _zz_cache_mru_3 = ways_3_metas_104_mru;
      end
      7'b1101001 : begin
        _zz_cache_tag_0 = ways_0_metas_105_tag;
        _zz_cache_hit_0 = ways_0_metas_105_vld;
        _zz_cache_mru_0 = ways_0_metas_105_mru;
        _zz_cache_tag_1 = ways_1_metas_105_tag;
        _zz_cache_hit_1 = ways_1_metas_105_vld;
        _zz_cache_mru_1 = ways_1_metas_105_mru;
        _zz_cache_tag_2 = ways_2_metas_105_tag;
        _zz_cache_hit_2 = ways_2_metas_105_vld;
        _zz_cache_mru_2 = ways_2_metas_105_mru;
        _zz_cache_tag_3 = ways_3_metas_105_tag;
        _zz_cache_hit_3 = ways_3_metas_105_vld;
        _zz_cache_mru_3 = ways_3_metas_105_mru;
      end
      7'b1101010 : begin
        _zz_cache_tag_0 = ways_0_metas_106_tag;
        _zz_cache_hit_0 = ways_0_metas_106_vld;
        _zz_cache_mru_0 = ways_0_metas_106_mru;
        _zz_cache_tag_1 = ways_1_metas_106_tag;
        _zz_cache_hit_1 = ways_1_metas_106_vld;
        _zz_cache_mru_1 = ways_1_metas_106_mru;
        _zz_cache_tag_2 = ways_2_metas_106_tag;
        _zz_cache_hit_2 = ways_2_metas_106_vld;
        _zz_cache_mru_2 = ways_2_metas_106_mru;
        _zz_cache_tag_3 = ways_3_metas_106_tag;
        _zz_cache_hit_3 = ways_3_metas_106_vld;
        _zz_cache_mru_3 = ways_3_metas_106_mru;
      end
      7'b1101011 : begin
        _zz_cache_tag_0 = ways_0_metas_107_tag;
        _zz_cache_hit_0 = ways_0_metas_107_vld;
        _zz_cache_mru_0 = ways_0_metas_107_mru;
        _zz_cache_tag_1 = ways_1_metas_107_tag;
        _zz_cache_hit_1 = ways_1_metas_107_vld;
        _zz_cache_mru_1 = ways_1_metas_107_mru;
        _zz_cache_tag_2 = ways_2_metas_107_tag;
        _zz_cache_hit_2 = ways_2_metas_107_vld;
        _zz_cache_mru_2 = ways_2_metas_107_mru;
        _zz_cache_tag_3 = ways_3_metas_107_tag;
        _zz_cache_hit_3 = ways_3_metas_107_vld;
        _zz_cache_mru_3 = ways_3_metas_107_mru;
      end
      7'b1101100 : begin
        _zz_cache_tag_0 = ways_0_metas_108_tag;
        _zz_cache_hit_0 = ways_0_metas_108_vld;
        _zz_cache_mru_0 = ways_0_metas_108_mru;
        _zz_cache_tag_1 = ways_1_metas_108_tag;
        _zz_cache_hit_1 = ways_1_metas_108_vld;
        _zz_cache_mru_1 = ways_1_metas_108_mru;
        _zz_cache_tag_2 = ways_2_metas_108_tag;
        _zz_cache_hit_2 = ways_2_metas_108_vld;
        _zz_cache_mru_2 = ways_2_metas_108_mru;
        _zz_cache_tag_3 = ways_3_metas_108_tag;
        _zz_cache_hit_3 = ways_3_metas_108_vld;
        _zz_cache_mru_3 = ways_3_metas_108_mru;
      end
      7'b1101101 : begin
        _zz_cache_tag_0 = ways_0_metas_109_tag;
        _zz_cache_hit_0 = ways_0_metas_109_vld;
        _zz_cache_mru_0 = ways_0_metas_109_mru;
        _zz_cache_tag_1 = ways_1_metas_109_tag;
        _zz_cache_hit_1 = ways_1_metas_109_vld;
        _zz_cache_mru_1 = ways_1_metas_109_mru;
        _zz_cache_tag_2 = ways_2_metas_109_tag;
        _zz_cache_hit_2 = ways_2_metas_109_vld;
        _zz_cache_mru_2 = ways_2_metas_109_mru;
        _zz_cache_tag_3 = ways_3_metas_109_tag;
        _zz_cache_hit_3 = ways_3_metas_109_vld;
        _zz_cache_mru_3 = ways_3_metas_109_mru;
      end
      7'b1101110 : begin
        _zz_cache_tag_0 = ways_0_metas_110_tag;
        _zz_cache_hit_0 = ways_0_metas_110_vld;
        _zz_cache_mru_0 = ways_0_metas_110_mru;
        _zz_cache_tag_1 = ways_1_metas_110_tag;
        _zz_cache_hit_1 = ways_1_metas_110_vld;
        _zz_cache_mru_1 = ways_1_metas_110_mru;
        _zz_cache_tag_2 = ways_2_metas_110_tag;
        _zz_cache_hit_2 = ways_2_metas_110_vld;
        _zz_cache_mru_2 = ways_2_metas_110_mru;
        _zz_cache_tag_3 = ways_3_metas_110_tag;
        _zz_cache_hit_3 = ways_3_metas_110_vld;
        _zz_cache_mru_3 = ways_3_metas_110_mru;
      end
      7'b1101111 : begin
        _zz_cache_tag_0 = ways_0_metas_111_tag;
        _zz_cache_hit_0 = ways_0_metas_111_vld;
        _zz_cache_mru_0 = ways_0_metas_111_mru;
        _zz_cache_tag_1 = ways_1_metas_111_tag;
        _zz_cache_hit_1 = ways_1_metas_111_vld;
        _zz_cache_mru_1 = ways_1_metas_111_mru;
        _zz_cache_tag_2 = ways_2_metas_111_tag;
        _zz_cache_hit_2 = ways_2_metas_111_vld;
        _zz_cache_mru_2 = ways_2_metas_111_mru;
        _zz_cache_tag_3 = ways_3_metas_111_tag;
        _zz_cache_hit_3 = ways_3_metas_111_vld;
        _zz_cache_mru_3 = ways_3_metas_111_mru;
      end
      7'b1110000 : begin
        _zz_cache_tag_0 = ways_0_metas_112_tag;
        _zz_cache_hit_0 = ways_0_metas_112_vld;
        _zz_cache_mru_0 = ways_0_metas_112_mru;
        _zz_cache_tag_1 = ways_1_metas_112_tag;
        _zz_cache_hit_1 = ways_1_metas_112_vld;
        _zz_cache_mru_1 = ways_1_metas_112_mru;
        _zz_cache_tag_2 = ways_2_metas_112_tag;
        _zz_cache_hit_2 = ways_2_metas_112_vld;
        _zz_cache_mru_2 = ways_2_metas_112_mru;
        _zz_cache_tag_3 = ways_3_metas_112_tag;
        _zz_cache_hit_3 = ways_3_metas_112_vld;
        _zz_cache_mru_3 = ways_3_metas_112_mru;
      end
      7'b1110001 : begin
        _zz_cache_tag_0 = ways_0_metas_113_tag;
        _zz_cache_hit_0 = ways_0_metas_113_vld;
        _zz_cache_mru_0 = ways_0_metas_113_mru;
        _zz_cache_tag_1 = ways_1_metas_113_tag;
        _zz_cache_hit_1 = ways_1_metas_113_vld;
        _zz_cache_mru_1 = ways_1_metas_113_mru;
        _zz_cache_tag_2 = ways_2_metas_113_tag;
        _zz_cache_hit_2 = ways_2_metas_113_vld;
        _zz_cache_mru_2 = ways_2_metas_113_mru;
        _zz_cache_tag_3 = ways_3_metas_113_tag;
        _zz_cache_hit_3 = ways_3_metas_113_vld;
        _zz_cache_mru_3 = ways_3_metas_113_mru;
      end
      7'b1110010 : begin
        _zz_cache_tag_0 = ways_0_metas_114_tag;
        _zz_cache_hit_0 = ways_0_metas_114_vld;
        _zz_cache_mru_0 = ways_0_metas_114_mru;
        _zz_cache_tag_1 = ways_1_metas_114_tag;
        _zz_cache_hit_1 = ways_1_metas_114_vld;
        _zz_cache_mru_1 = ways_1_metas_114_mru;
        _zz_cache_tag_2 = ways_2_metas_114_tag;
        _zz_cache_hit_2 = ways_2_metas_114_vld;
        _zz_cache_mru_2 = ways_2_metas_114_mru;
        _zz_cache_tag_3 = ways_3_metas_114_tag;
        _zz_cache_hit_3 = ways_3_metas_114_vld;
        _zz_cache_mru_3 = ways_3_metas_114_mru;
      end
      7'b1110011 : begin
        _zz_cache_tag_0 = ways_0_metas_115_tag;
        _zz_cache_hit_0 = ways_0_metas_115_vld;
        _zz_cache_mru_0 = ways_0_metas_115_mru;
        _zz_cache_tag_1 = ways_1_metas_115_tag;
        _zz_cache_hit_1 = ways_1_metas_115_vld;
        _zz_cache_mru_1 = ways_1_metas_115_mru;
        _zz_cache_tag_2 = ways_2_metas_115_tag;
        _zz_cache_hit_2 = ways_2_metas_115_vld;
        _zz_cache_mru_2 = ways_2_metas_115_mru;
        _zz_cache_tag_3 = ways_3_metas_115_tag;
        _zz_cache_hit_3 = ways_3_metas_115_vld;
        _zz_cache_mru_3 = ways_3_metas_115_mru;
      end
      7'b1110100 : begin
        _zz_cache_tag_0 = ways_0_metas_116_tag;
        _zz_cache_hit_0 = ways_0_metas_116_vld;
        _zz_cache_mru_0 = ways_0_metas_116_mru;
        _zz_cache_tag_1 = ways_1_metas_116_tag;
        _zz_cache_hit_1 = ways_1_metas_116_vld;
        _zz_cache_mru_1 = ways_1_metas_116_mru;
        _zz_cache_tag_2 = ways_2_metas_116_tag;
        _zz_cache_hit_2 = ways_2_metas_116_vld;
        _zz_cache_mru_2 = ways_2_metas_116_mru;
        _zz_cache_tag_3 = ways_3_metas_116_tag;
        _zz_cache_hit_3 = ways_3_metas_116_vld;
        _zz_cache_mru_3 = ways_3_metas_116_mru;
      end
      7'b1110101 : begin
        _zz_cache_tag_0 = ways_0_metas_117_tag;
        _zz_cache_hit_0 = ways_0_metas_117_vld;
        _zz_cache_mru_0 = ways_0_metas_117_mru;
        _zz_cache_tag_1 = ways_1_metas_117_tag;
        _zz_cache_hit_1 = ways_1_metas_117_vld;
        _zz_cache_mru_1 = ways_1_metas_117_mru;
        _zz_cache_tag_2 = ways_2_metas_117_tag;
        _zz_cache_hit_2 = ways_2_metas_117_vld;
        _zz_cache_mru_2 = ways_2_metas_117_mru;
        _zz_cache_tag_3 = ways_3_metas_117_tag;
        _zz_cache_hit_3 = ways_3_metas_117_vld;
        _zz_cache_mru_3 = ways_3_metas_117_mru;
      end
      7'b1110110 : begin
        _zz_cache_tag_0 = ways_0_metas_118_tag;
        _zz_cache_hit_0 = ways_0_metas_118_vld;
        _zz_cache_mru_0 = ways_0_metas_118_mru;
        _zz_cache_tag_1 = ways_1_metas_118_tag;
        _zz_cache_hit_1 = ways_1_metas_118_vld;
        _zz_cache_mru_1 = ways_1_metas_118_mru;
        _zz_cache_tag_2 = ways_2_metas_118_tag;
        _zz_cache_hit_2 = ways_2_metas_118_vld;
        _zz_cache_mru_2 = ways_2_metas_118_mru;
        _zz_cache_tag_3 = ways_3_metas_118_tag;
        _zz_cache_hit_3 = ways_3_metas_118_vld;
        _zz_cache_mru_3 = ways_3_metas_118_mru;
      end
      7'b1110111 : begin
        _zz_cache_tag_0 = ways_0_metas_119_tag;
        _zz_cache_hit_0 = ways_0_metas_119_vld;
        _zz_cache_mru_0 = ways_0_metas_119_mru;
        _zz_cache_tag_1 = ways_1_metas_119_tag;
        _zz_cache_hit_1 = ways_1_metas_119_vld;
        _zz_cache_mru_1 = ways_1_metas_119_mru;
        _zz_cache_tag_2 = ways_2_metas_119_tag;
        _zz_cache_hit_2 = ways_2_metas_119_vld;
        _zz_cache_mru_2 = ways_2_metas_119_mru;
        _zz_cache_tag_3 = ways_3_metas_119_tag;
        _zz_cache_hit_3 = ways_3_metas_119_vld;
        _zz_cache_mru_3 = ways_3_metas_119_mru;
      end
      7'b1111000 : begin
        _zz_cache_tag_0 = ways_0_metas_120_tag;
        _zz_cache_hit_0 = ways_0_metas_120_vld;
        _zz_cache_mru_0 = ways_0_metas_120_mru;
        _zz_cache_tag_1 = ways_1_metas_120_tag;
        _zz_cache_hit_1 = ways_1_metas_120_vld;
        _zz_cache_mru_1 = ways_1_metas_120_mru;
        _zz_cache_tag_2 = ways_2_metas_120_tag;
        _zz_cache_hit_2 = ways_2_metas_120_vld;
        _zz_cache_mru_2 = ways_2_metas_120_mru;
        _zz_cache_tag_3 = ways_3_metas_120_tag;
        _zz_cache_hit_3 = ways_3_metas_120_vld;
        _zz_cache_mru_3 = ways_3_metas_120_mru;
      end
      7'b1111001 : begin
        _zz_cache_tag_0 = ways_0_metas_121_tag;
        _zz_cache_hit_0 = ways_0_metas_121_vld;
        _zz_cache_mru_0 = ways_0_metas_121_mru;
        _zz_cache_tag_1 = ways_1_metas_121_tag;
        _zz_cache_hit_1 = ways_1_metas_121_vld;
        _zz_cache_mru_1 = ways_1_metas_121_mru;
        _zz_cache_tag_2 = ways_2_metas_121_tag;
        _zz_cache_hit_2 = ways_2_metas_121_vld;
        _zz_cache_mru_2 = ways_2_metas_121_mru;
        _zz_cache_tag_3 = ways_3_metas_121_tag;
        _zz_cache_hit_3 = ways_3_metas_121_vld;
        _zz_cache_mru_3 = ways_3_metas_121_mru;
      end
      7'b1111010 : begin
        _zz_cache_tag_0 = ways_0_metas_122_tag;
        _zz_cache_hit_0 = ways_0_metas_122_vld;
        _zz_cache_mru_0 = ways_0_metas_122_mru;
        _zz_cache_tag_1 = ways_1_metas_122_tag;
        _zz_cache_hit_1 = ways_1_metas_122_vld;
        _zz_cache_mru_1 = ways_1_metas_122_mru;
        _zz_cache_tag_2 = ways_2_metas_122_tag;
        _zz_cache_hit_2 = ways_2_metas_122_vld;
        _zz_cache_mru_2 = ways_2_metas_122_mru;
        _zz_cache_tag_3 = ways_3_metas_122_tag;
        _zz_cache_hit_3 = ways_3_metas_122_vld;
        _zz_cache_mru_3 = ways_3_metas_122_mru;
      end
      7'b1111011 : begin
        _zz_cache_tag_0 = ways_0_metas_123_tag;
        _zz_cache_hit_0 = ways_0_metas_123_vld;
        _zz_cache_mru_0 = ways_0_metas_123_mru;
        _zz_cache_tag_1 = ways_1_metas_123_tag;
        _zz_cache_hit_1 = ways_1_metas_123_vld;
        _zz_cache_mru_1 = ways_1_metas_123_mru;
        _zz_cache_tag_2 = ways_2_metas_123_tag;
        _zz_cache_hit_2 = ways_2_metas_123_vld;
        _zz_cache_mru_2 = ways_2_metas_123_mru;
        _zz_cache_tag_3 = ways_3_metas_123_tag;
        _zz_cache_hit_3 = ways_3_metas_123_vld;
        _zz_cache_mru_3 = ways_3_metas_123_mru;
      end
      7'b1111100 : begin
        _zz_cache_tag_0 = ways_0_metas_124_tag;
        _zz_cache_hit_0 = ways_0_metas_124_vld;
        _zz_cache_mru_0 = ways_0_metas_124_mru;
        _zz_cache_tag_1 = ways_1_metas_124_tag;
        _zz_cache_hit_1 = ways_1_metas_124_vld;
        _zz_cache_mru_1 = ways_1_metas_124_mru;
        _zz_cache_tag_2 = ways_2_metas_124_tag;
        _zz_cache_hit_2 = ways_2_metas_124_vld;
        _zz_cache_mru_2 = ways_2_metas_124_mru;
        _zz_cache_tag_3 = ways_3_metas_124_tag;
        _zz_cache_hit_3 = ways_3_metas_124_vld;
        _zz_cache_mru_3 = ways_3_metas_124_mru;
      end
      7'b1111101 : begin
        _zz_cache_tag_0 = ways_0_metas_125_tag;
        _zz_cache_hit_0 = ways_0_metas_125_vld;
        _zz_cache_mru_0 = ways_0_metas_125_mru;
        _zz_cache_tag_1 = ways_1_metas_125_tag;
        _zz_cache_hit_1 = ways_1_metas_125_vld;
        _zz_cache_mru_1 = ways_1_metas_125_mru;
        _zz_cache_tag_2 = ways_2_metas_125_tag;
        _zz_cache_hit_2 = ways_2_metas_125_vld;
        _zz_cache_mru_2 = ways_2_metas_125_mru;
        _zz_cache_tag_3 = ways_3_metas_125_tag;
        _zz_cache_hit_3 = ways_3_metas_125_vld;
        _zz_cache_mru_3 = ways_3_metas_125_mru;
      end
      7'b1111110 : begin
        _zz_cache_tag_0 = ways_0_metas_126_tag;
        _zz_cache_hit_0 = ways_0_metas_126_vld;
        _zz_cache_mru_0 = ways_0_metas_126_mru;
        _zz_cache_tag_1 = ways_1_metas_126_tag;
        _zz_cache_hit_1 = ways_1_metas_126_vld;
        _zz_cache_mru_1 = ways_1_metas_126_mru;
        _zz_cache_tag_2 = ways_2_metas_126_tag;
        _zz_cache_hit_2 = ways_2_metas_126_vld;
        _zz_cache_mru_2 = ways_2_metas_126_mru;
        _zz_cache_tag_3 = ways_3_metas_126_tag;
        _zz_cache_hit_3 = ways_3_metas_126_vld;
        _zz_cache_mru_3 = ways_3_metas_126_mru;
      end
      default : begin
        _zz_cache_tag_0 = ways_0_metas_127_tag;
        _zz_cache_hit_0 = ways_0_metas_127_vld;
        _zz_cache_mru_0 = ways_0_metas_127_mru;
        _zz_cache_tag_1 = ways_1_metas_127_tag;
        _zz_cache_hit_1 = ways_1_metas_127_vld;
        _zz_cache_mru_1 = ways_1_metas_127_mru;
        _zz_cache_tag_2 = ways_2_metas_127_tag;
        _zz_cache_hit_2 = ways_2_metas_127_vld;
        _zz_cache_mru_2 = ways_2_metas_127_mru;
        _zz_cache_tag_3 = ways_3_metas_127_tag;
        _zz_cache_hit_3 = ways_3_metas_127_vld;
        _zz_cache_mru_3 = ways_3_metas_127_mru;
      end
    endcase
  end

  always @(*) begin
    case(cpu_set_d1)
      7'b0000000 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_0_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_0_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_0_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_0_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_0_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_0_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_0_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_0_mru;
      end
      7'b0000001 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_1_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_1_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_1_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_1_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_1_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_1_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_1_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_1_mru;
      end
      7'b0000010 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_2_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_2_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_2_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_2_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_2_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_2_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_2_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_2_mru;
      end
      7'b0000011 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_3_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_3_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_3_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_3_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_3_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_3_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_3_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_3_mru;
      end
      7'b0000100 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_4_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_4_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_4_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_4_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_4_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_4_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_4_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_4_mru;
      end
      7'b0000101 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_5_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_5_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_5_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_5_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_5_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_5_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_5_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_5_mru;
      end
      7'b0000110 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_6_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_6_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_6_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_6_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_6_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_6_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_6_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_6_mru;
      end
      7'b0000111 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_7_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_7_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_7_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_7_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_7_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_7_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_7_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_7_mru;
      end
      7'b0001000 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_8_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_8_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_8_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_8_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_8_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_8_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_8_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_8_mru;
      end
      7'b0001001 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_9_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_9_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_9_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_9_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_9_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_9_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_9_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_9_mru;
      end
      7'b0001010 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_10_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_10_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_10_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_10_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_10_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_10_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_10_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_10_mru;
      end
      7'b0001011 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_11_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_11_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_11_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_11_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_11_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_11_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_11_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_11_mru;
      end
      7'b0001100 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_12_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_12_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_12_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_12_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_12_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_12_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_12_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_12_mru;
      end
      7'b0001101 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_13_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_13_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_13_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_13_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_13_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_13_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_13_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_13_mru;
      end
      7'b0001110 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_14_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_14_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_14_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_14_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_14_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_14_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_14_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_14_mru;
      end
      7'b0001111 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_15_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_15_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_15_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_15_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_15_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_15_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_15_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_15_mru;
      end
      7'b0010000 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_16_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_16_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_16_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_16_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_16_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_16_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_16_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_16_mru;
      end
      7'b0010001 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_17_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_17_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_17_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_17_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_17_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_17_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_17_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_17_mru;
      end
      7'b0010010 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_18_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_18_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_18_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_18_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_18_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_18_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_18_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_18_mru;
      end
      7'b0010011 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_19_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_19_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_19_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_19_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_19_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_19_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_19_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_19_mru;
      end
      7'b0010100 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_20_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_20_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_20_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_20_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_20_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_20_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_20_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_20_mru;
      end
      7'b0010101 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_21_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_21_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_21_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_21_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_21_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_21_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_21_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_21_mru;
      end
      7'b0010110 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_22_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_22_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_22_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_22_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_22_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_22_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_22_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_22_mru;
      end
      7'b0010111 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_23_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_23_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_23_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_23_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_23_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_23_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_23_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_23_mru;
      end
      7'b0011000 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_24_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_24_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_24_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_24_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_24_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_24_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_24_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_24_mru;
      end
      7'b0011001 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_25_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_25_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_25_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_25_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_25_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_25_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_25_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_25_mru;
      end
      7'b0011010 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_26_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_26_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_26_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_26_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_26_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_26_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_26_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_26_mru;
      end
      7'b0011011 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_27_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_27_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_27_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_27_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_27_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_27_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_27_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_27_mru;
      end
      7'b0011100 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_28_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_28_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_28_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_28_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_28_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_28_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_28_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_28_mru;
      end
      7'b0011101 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_29_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_29_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_29_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_29_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_29_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_29_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_29_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_29_mru;
      end
      7'b0011110 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_30_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_30_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_30_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_30_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_30_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_30_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_30_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_30_mru;
      end
      7'b0011111 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_31_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_31_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_31_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_31_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_31_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_31_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_31_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_31_mru;
      end
      7'b0100000 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_32_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_32_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_32_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_32_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_32_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_32_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_32_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_32_mru;
      end
      7'b0100001 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_33_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_33_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_33_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_33_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_33_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_33_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_33_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_33_mru;
      end
      7'b0100010 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_34_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_34_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_34_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_34_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_34_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_34_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_34_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_34_mru;
      end
      7'b0100011 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_35_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_35_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_35_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_35_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_35_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_35_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_35_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_35_mru;
      end
      7'b0100100 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_36_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_36_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_36_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_36_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_36_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_36_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_36_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_36_mru;
      end
      7'b0100101 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_37_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_37_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_37_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_37_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_37_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_37_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_37_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_37_mru;
      end
      7'b0100110 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_38_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_38_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_38_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_38_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_38_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_38_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_38_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_38_mru;
      end
      7'b0100111 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_39_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_39_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_39_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_39_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_39_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_39_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_39_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_39_mru;
      end
      7'b0101000 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_40_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_40_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_40_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_40_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_40_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_40_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_40_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_40_mru;
      end
      7'b0101001 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_41_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_41_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_41_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_41_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_41_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_41_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_41_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_41_mru;
      end
      7'b0101010 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_42_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_42_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_42_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_42_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_42_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_42_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_42_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_42_mru;
      end
      7'b0101011 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_43_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_43_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_43_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_43_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_43_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_43_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_43_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_43_mru;
      end
      7'b0101100 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_44_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_44_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_44_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_44_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_44_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_44_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_44_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_44_mru;
      end
      7'b0101101 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_45_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_45_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_45_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_45_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_45_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_45_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_45_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_45_mru;
      end
      7'b0101110 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_46_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_46_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_46_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_46_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_46_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_46_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_46_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_46_mru;
      end
      7'b0101111 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_47_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_47_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_47_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_47_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_47_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_47_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_47_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_47_mru;
      end
      7'b0110000 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_48_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_48_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_48_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_48_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_48_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_48_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_48_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_48_mru;
      end
      7'b0110001 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_49_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_49_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_49_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_49_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_49_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_49_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_49_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_49_mru;
      end
      7'b0110010 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_50_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_50_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_50_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_50_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_50_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_50_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_50_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_50_mru;
      end
      7'b0110011 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_51_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_51_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_51_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_51_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_51_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_51_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_51_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_51_mru;
      end
      7'b0110100 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_52_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_52_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_52_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_52_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_52_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_52_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_52_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_52_mru;
      end
      7'b0110101 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_53_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_53_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_53_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_53_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_53_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_53_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_53_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_53_mru;
      end
      7'b0110110 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_54_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_54_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_54_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_54_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_54_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_54_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_54_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_54_mru;
      end
      7'b0110111 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_55_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_55_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_55_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_55_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_55_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_55_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_55_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_55_mru;
      end
      7'b0111000 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_56_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_56_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_56_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_56_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_56_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_56_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_56_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_56_mru;
      end
      7'b0111001 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_57_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_57_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_57_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_57_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_57_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_57_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_57_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_57_mru;
      end
      7'b0111010 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_58_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_58_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_58_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_58_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_58_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_58_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_58_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_58_mru;
      end
      7'b0111011 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_59_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_59_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_59_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_59_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_59_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_59_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_59_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_59_mru;
      end
      7'b0111100 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_60_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_60_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_60_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_60_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_60_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_60_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_60_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_60_mru;
      end
      7'b0111101 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_61_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_61_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_61_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_61_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_61_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_61_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_61_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_61_mru;
      end
      7'b0111110 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_62_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_62_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_62_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_62_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_62_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_62_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_62_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_62_mru;
      end
      7'b0111111 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_63_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_63_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_63_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_63_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_63_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_63_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_63_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_63_mru;
      end
      7'b1000000 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_64_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_64_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_64_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_64_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_64_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_64_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_64_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_64_mru;
      end
      7'b1000001 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_65_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_65_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_65_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_65_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_65_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_65_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_65_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_65_mru;
      end
      7'b1000010 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_66_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_66_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_66_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_66_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_66_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_66_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_66_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_66_mru;
      end
      7'b1000011 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_67_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_67_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_67_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_67_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_67_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_67_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_67_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_67_mru;
      end
      7'b1000100 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_68_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_68_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_68_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_68_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_68_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_68_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_68_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_68_mru;
      end
      7'b1000101 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_69_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_69_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_69_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_69_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_69_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_69_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_69_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_69_mru;
      end
      7'b1000110 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_70_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_70_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_70_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_70_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_70_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_70_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_70_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_70_mru;
      end
      7'b1000111 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_71_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_71_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_71_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_71_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_71_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_71_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_71_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_71_mru;
      end
      7'b1001000 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_72_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_72_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_72_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_72_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_72_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_72_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_72_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_72_mru;
      end
      7'b1001001 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_73_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_73_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_73_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_73_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_73_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_73_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_73_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_73_mru;
      end
      7'b1001010 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_74_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_74_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_74_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_74_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_74_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_74_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_74_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_74_mru;
      end
      7'b1001011 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_75_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_75_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_75_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_75_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_75_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_75_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_75_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_75_mru;
      end
      7'b1001100 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_76_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_76_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_76_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_76_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_76_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_76_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_76_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_76_mru;
      end
      7'b1001101 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_77_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_77_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_77_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_77_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_77_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_77_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_77_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_77_mru;
      end
      7'b1001110 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_78_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_78_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_78_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_78_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_78_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_78_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_78_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_78_mru;
      end
      7'b1001111 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_79_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_79_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_79_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_79_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_79_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_79_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_79_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_79_mru;
      end
      7'b1010000 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_80_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_80_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_80_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_80_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_80_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_80_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_80_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_80_mru;
      end
      7'b1010001 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_81_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_81_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_81_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_81_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_81_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_81_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_81_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_81_mru;
      end
      7'b1010010 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_82_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_82_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_82_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_82_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_82_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_82_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_82_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_82_mru;
      end
      7'b1010011 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_83_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_83_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_83_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_83_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_83_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_83_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_83_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_83_mru;
      end
      7'b1010100 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_84_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_84_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_84_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_84_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_84_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_84_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_84_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_84_mru;
      end
      7'b1010101 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_85_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_85_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_85_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_85_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_85_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_85_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_85_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_85_mru;
      end
      7'b1010110 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_86_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_86_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_86_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_86_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_86_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_86_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_86_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_86_mru;
      end
      7'b1010111 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_87_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_87_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_87_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_87_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_87_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_87_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_87_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_87_mru;
      end
      7'b1011000 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_88_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_88_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_88_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_88_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_88_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_88_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_88_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_88_mru;
      end
      7'b1011001 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_89_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_89_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_89_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_89_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_89_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_89_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_89_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_89_mru;
      end
      7'b1011010 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_90_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_90_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_90_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_90_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_90_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_90_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_90_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_90_mru;
      end
      7'b1011011 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_91_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_91_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_91_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_91_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_91_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_91_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_91_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_91_mru;
      end
      7'b1011100 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_92_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_92_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_92_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_92_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_92_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_92_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_92_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_92_mru;
      end
      7'b1011101 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_93_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_93_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_93_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_93_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_93_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_93_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_93_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_93_mru;
      end
      7'b1011110 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_94_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_94_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_94_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_94_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_94_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_94_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_94_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_94_mru;
      end
      7'b1011111 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_95_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_95_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_95_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_95_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_95_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_95_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_95_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_95_mru;
      end
      7'b1100000 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_96_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_96_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_96_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_96_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_96_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_96_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_96_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_96_mru;
      end
      7'b1100001 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_97_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_97_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_97_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_97_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_97_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_97_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_97_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_97_mru;
      end
      7'b1100010 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_98_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_98_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_98_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_98_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_98_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_98_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_98_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_98_mru;
      end
      7'b1100011 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_99_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_99_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_99_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_99_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_99_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_99_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_99_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_99_mru;
      end
      7'b1100100 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_100_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_100_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_100_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_100_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_100_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_100_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_100_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_100_mru;
      end
      7'b1100101 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_101_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_101_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_101_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_101_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_101_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_101_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_101_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_101_mru;
      end
      7'b1100110 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_102_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_102_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_102_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_102_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_102_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_102_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_102_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_102_mru;
      end
      7'b1100111 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_103_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_103_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_103_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_103_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_103_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_103_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_103_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_103_mru;
      end
      7'b1101000 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_104_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_104_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_104_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_104_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_104_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_104_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_104_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_104_mru;
      end
      7'b1101001 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_105_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_105_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_105_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_105_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_105_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_105_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_105_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_105_mru;
      end
      7'b1101010 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_106_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_106_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_106_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_106_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_106_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_106_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_106_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_106_mru;
      end
      7'b1101011 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_107_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_107_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_107_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_107_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_107_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_107_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_107_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_107_mru;
      end
      7'b1101100 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_108_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_108_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_108_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_108_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_108_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_108_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_108_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_108_mru;
      end
      7'b1101101 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_109_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_109_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_109_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_109_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_109_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_109_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_109_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_109_mru;
      end
      7'b1101110 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_110_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_110_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_110_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_110_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_110_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_110_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_110_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_110_mru;
      end
      7'b1101111 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_111_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_111_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_111_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_111_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_111_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_111_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_111_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_111_mru;
      end
      7'b1110000 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_112_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_112_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_112_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_112_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_112_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_112_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_112_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_112_mru;
      end
      7'b1110001 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_113_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_113_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_113_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_113_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_113_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_113_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_113_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_113_mru;
      end
      7'b1110010 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_114_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_114_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_114_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_114_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_114_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_114_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_114_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_114_mru;
      end
      7'b1110011 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_115_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_115_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_115_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_115_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_115_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_115_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_115_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_115_mru;
      end
      7'b1110100 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_116_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_116_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_116_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_116_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_116_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_116_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_116_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_116_mru;
      end
      7'b1110101 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_117_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_117_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_117_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_117_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_117_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_117_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_117_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_117_mru;
      end
      7'b1110110 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_118_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_118_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_118_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_118_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_118_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_118_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_118_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_118_mru;
      end
      7'b1110111 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_119_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_119_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_119_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_119_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_119_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_119_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_119_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_119_mru;
      end
      7'b1111000 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_120_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_120_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_120_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_120_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_120_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_120_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_120_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_120_mru;
      end
      7'b1111001 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_121_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_121_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_121_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_121_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_121_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_121_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_121_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_121_mru;
      end
      7'b1111010 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_122_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_122_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_122_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_122_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_122_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_122_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_122_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_122_mru;
      end
      7'b1111011 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_123_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_123_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_123_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_123_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_123_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_123_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_123_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_123_mru;
      end
      7'b1111100 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_124_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_124_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_124_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_124_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_124_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_124_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_124_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_124_mru;
      end
      7'b1111101 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_125_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_125_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_125_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_125_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_125_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_125_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_125_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_125_mru;
      end
      7'b1111110 : begin
        _zz_cache_invld_d1_0 = ways_0_metas_126_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_126_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_126_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_126_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_126_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_126_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_126_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_126_mru;
      end
      default : begin
        _zz_cache_invld_d1_0 = ways_0_metas_127_vld;
        _zz_cache_lru_d1_0 = ways_0_metas_127_mru;
        _zz_cache_invld_d1_1 = ways_1_metas_127_vld;
        _zz_cache_lru_d1_1 = ways_1_metas_127_mru;
        _zz_cache_invld_d1_2 = ways_2_metas_127_vld;
        _zz_cache_lru_d1_2 = ways_2_metas_127_mru;
        _zz_cache_invld_d1_3 = ways_3_metas_127_vld;
        _zz_cache_lru_d1_3 = ways_3_metas_127_mru;
      end
    endcase
  end

  always @(*) begin
    case(hit_id_d1)
      2'b00 : begin
        _zz__zz_cpu_rsp_payload_data = sram_banks_data_0;
        _zz_cpu_rsp_valid = sram_banks_valid_0;
      end
      2'b01 : begin
        _zz__zz_cpu_rsp_payload_data = sram_banks_data_1;
        _zz_cpu_rsp_valid = sram_banks_valid_1;
      end
      2'b10 : begin
        _zz__zz_cpu_rsp_payload_data = sram_banks_data_2;
        _zz_cpu_rsp_valid = sram_banks_valid_2;
      end
      default : begin
        _zz__zz_cpu_rsp_payload_data = sram_banks_data_3;
        _zz_cpu_rsp_valid = sram_banks_valid_3;
      end
    endcase
  end

  always @(*) begin
    case(evict_id_miss)
      2'b00 : begin
        _zz__zz_cpu_rsp_payload_data_1 = sram_banks_data_0;
        _zz_cpu_rsp_valid_1 = sram_banks_valid_0;
      end
      2'b01 : begin
        _zz__zz_cpu_rsp_payload_data_1 = sram_banks_data_1;
        _zz_cpu_rsp_valid_1 = sram_banks_valid_1;
      end
      2'b10 : begin
        _zz__zz_cpu_rsp_payload_data_1 = sram_banks_data_2;
        _zz_cpu_rsp_valid_1 = sram_banks_valid_2;
      end
      default : begin
        _zz__zz_cpu_rsp_payload_data_1 = sram_banks_data_3;
        _zz_cpu_rsp_valid_1 = sram_banks_valid_3;
      end
    endcase
  end

  always @(*) begin
    case(cpu_bank_index_d1)
      4'b0000 : begin
        _zz_cpu_rsp_payload_data_2 = _zz_cpu_rsp_payload_data[31 : 0];
        _zz_cpu_rsp_payload_data_3 = _zz_cpu_rsp_payload_data_1[31 : 0];
      end
      4'b0001 : begin
        _zz_cpu_rsp_payload_data_2 = _zz_cpu_rsp_payload_data[63 : 32];
        _zz_cpu_rsp_payload_data_3 = _zz_cpu_rsp_payload_data_1[63 : 32];
      end
      4'b0010 : begin
        _zz_cpu_rsp_payload_data_2 = _zz_cpu_rsp_payload_data[95 : 64];
        _zz_cpu_rsp_payload_data_3 = _zz_cpu_rsp_payload_data_1[95 : 64];
      end
      4'b0011 : begin
        _zz_cpu_rsp_payload_data_2 = _zz_cpu_rsp_payload_data[127 : 96];
        _zz_cpu_rsp_payload_data_3 = _zz_cpu_rsp_payload_data_1[127 : 96];
      end
      4'b0100 : begin
        _zz_cpu_rsp_payload_data_2 = _zz_cpu_rsp_payload_data[159 : 128];
        _zz_cpu_rsp_payload_data_3 = _zz_cpu_rsp_payload_data_1[159 : 128];
      end
      4'b0101 : begin
        _zz_cpu_rsp_payload_data_2 = _zz_cpu_rsp_payload_data[191 : 160];
        _zz_cpu_rsp_payload_data_3 = _zz_cpu_rsp_payload_data_1[191 : 160];
      end
      4'b0110 : begin
        _zz_cpu_rsp_payload_data_2 = _zz_cpu_rsp_payload_data[223 : 192];
        _zz_cpu_rsp_payload_data_3 = _zz_cpu_rsp_payload_data_1[223 : 192];
      end
      4'b0111 : begin
        _zz_cpu_rsp_payload_data_2 = _zz_cpu_rsp_payload_data[255 : 224];
        _zz_cpu_rsp_payload_data_3 = _zz_cpu_rsp_payload_data_1[255 : 224];
      end
      4'b1000 : begin
        _zz_cpu_rsp_payload_data_2 = _zz_cpu_rsp_payload_data[287 : 256];
        _zz_cpu_rsp_payload_data_3 = _zz_cpu_rsp_payload_data_1[287 : 256];
      end
      4'b1001 : begin
        _zz_cpu_rsp_payload_data_2 = _zz_cpu_rsp_payload_data[319 : 288];
        _zz_cpu_rsp_payload_data_3 = _zz_cpu_rsp_payload_data_1[319 : 288];
      end
      4'b1010 : begin
        _zz_cpu_rsp_payload_data_2 = _zz_cpu_rsp_payload_data[351 : 320];
        _zz_cpu_rsp_payload_data_3 = _zz_cpu_rsp_payload_data_1[351 : 320];
      end
      4'b1011 : begin
        _zz_cpu_rsp_payload_data_2 = _zz_cpu_rsp_payload_data[383 : 352];
        _zz_cpu_rsp_payload_data_3 = _zz_cpu_rsp_payload_data_1[383 : 352];
      end
      4'b1100 : begin
        _zz_cpu_rsp_payload_data_2 = _zz_cpu_rsp_payload_data[415 : 384];
        _zz_cpu_rsp_payload_data_3 = _zz_cpu_rsp_payload_data_1[415 : 384];
      end
      4'b1101 : begin
        _zz_cpu_rsp_payload_data_2 = _zz_cpu_rsp_payload_data[447 : 416];
        _zz_cpu_rsp_payload_data_3 = _zz_cpu_rsp_payload_data_1[447 : 416];
      end
      4'b1110 : begin
        _zz_cpu_rsp_payload_data_2 = _zz_cpu_rsp_payload_data[479 : 448];
        _zz_cpu_rsp_payload_data_3 = _zz_cpu_rsp_payload_data_1[479 : 448];
      end
      default : begin
        _zz_cpu_rsp_payload_data_2 = _zz_cpu_rsp_payload_data[511 : 480];
        _zz_cpu_rsp_payload_data_3 = _zz_cpu_rsp_payload_data_1[511 : 480];
      end
    endcase
  end

  assign mru_full = (&{cache_mru_3,{cache_mru_2,{cache_mru_1,cache_mru_0}}});
  assign cpu_cmd_fire = (cpu_cmd_valid && cpu_cmd_ready);
  assign is_hit = ((|{cache_hit_3,{cache_hit_2,{cache_hit_1,cache_hit_0}}}) && cpu_cmd_fire);
  assign cpu_cmd_fire_1 = (cpu_cmd_valid && cpu_cmd_ready);
  assign is_miss = ((! (|{cache_hit_3,{cache_hit_2,{cache_hit_1,cache_hit_0}}})) && cpu_cmd_fire_1);
  assign is_diff = (! (|{cache_victim_3,{cache_victim_2,{cache_victim_1,cache_victim_0}}}));
  always @(*) begin
    flush_cnt_willIncrement = 1'b0;
    if(!when_ICache_l142) begin
      if(flush_busy) begin
        flush_cnt_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    flush_cnt_willClear = 1'b0;
    if(when_ICache_l142) begin
      flush_cnt_willClear = 1'b1;
    end
  end

  assign flush_cnt_willOverflowIfInc = (flush_cnt_value == 7'h7f);
  assign flush_cnt_willOverflow = (flush_cnt_willOverflowIfInc && flush_cnt_willIncrement);
  always @(*) begin
    flush_cnt_valueNext = (flush_cnt_value + _zz_flush_cnt_valueNext);
    if(flush_cnt_willClear) begin
      flush_cnt_valueNext = 7'h0;
    end
  end

  assign flush_done = (flush_busy && (flush_cnt_value == 7'h7f));
  assign cpu_tag = cpu_cmd_payload_addr[63 : 13];
  assign cpu_set = cpu_cmd_payload_addr[12 : 6];
  assign cpu_bank_addr = cpu_cmd_payload_addr[12 : 6];
  assign cpu_bank_index = cpu_cmd_payload_addr[5 : 2];
  assign cpu_cmd_fire_2 = (cpu_cmd_valid && cpu_cmd_ready);
  assign cpu_set_d1 = cpu_addr_d1[12 : 6];
  assign cpu_tag_d1 = cpu_addr_d1[63 : 13];
  assign cpu_bank_addr_d1 = cpu_addr_d1[12 : 6];
  assign cpu_bank_index_d1 = cpu_addr_d1[5 : 2];
  always @(*) begin
    next_level_data_cnt_willIncrement = 1'b0;
    if(!is_miss) begin
      if(!next_level_done) begin
        if(next_level_rsp_valid) begin
          next_level_data_cnt_willIncrement = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    next_level_data_cnt_willClear = 1'b0;
    if(is_miss) begin
      next_level_data_cnt_willClear = 1'b1;
    end else begin
      if(next_level_done) begin
        next_level_data_cnt_willClear = 1'b1;
      end
    end
  end

  assign next_level_data_cnt_willOverflowIfInc = (next_level_data_cnt_value == 3'b111);
  assign next_level_data_cnt_willOverflow = (next_level_data_cnt_willOverflowIfInc && next_level_data_cnt_willIncrement);
  always @(*) begin
    next_level_data_cnt_valueNext = (next_level_data_cnt_value + _zz_next_level_data_cnt_valueNext);
    if(next_level_data_cnt_willClear) begin
      next_level_data_cnt_valueNext = 3'b000;
    end
  end

  assign next_level_bank_addr = cpu_addr_d1[12 : 6];
  assign next_level_cmd_fire = (next_level_cmd_valid && next_level_cmd_ready);
  assign when_ICache_l142 = (flush_busy && (flush_cnt_value == 7'h7f));
  assign _zz_cache_hit_gnt_0 = 4'b0001;
  assign _zz_cache_hit_gnt_0_1 = {cache_hit_3,{cache_hit_2,{cache_hit_1,cache_hit_0}}};
  assign _zz_cache_hit_gnt_0_2 = {_zz_cache_hit_gnt_0_1,_zz_cache_hit_gnt_0_1};
  assign _zz_cache_hit_gnt_0_3 = (_zz_cache_hit_gnt_0_2 & (~ _zz__zz_cache_hit_gnt_0_3));
  assign _zz_cache_hit_gnt_0_4 = (_zz_cache_hit_gnt_0_3[7 : 4] | _zz_cache_hit_gnt_0_3[3 : 0]);
  assign cache_hit_gnt_0 = _zz_cache_hit_gnt_0_4[0];
  assign cache_hit_gnt_1 = _zz_cache_hit_gnt_0_4[1];
  assign cache_hit_gnt_2 = _zz_cache_hit_gnt_0_4[2];
  assign cache_hit_gnt_3 = _zz_cache_hit_gnt_0_4[3];
  assign _zz_cache_invld_gnt_0 = 4'b0001;
  assign _zz_cache_invld_gnt_0_1 = {cache_invld_d1_3,{cache_invld_d1_2,{cache_invld_d1_1,cache_invld_d1_0}}};
  assign _zz_cache_invld_gnt_0_2 = {_zz_cache_invld_gnt_0_1,_zz_cache_invld_gnt_0_1};
  assign _zz_cache_invld_gnt_0_3 = (_zz_cache_invld_gnt_0_2 & (~ _zz__zz_cache_invld_gnt_0_3));
  assign _zz_cache_invld_gnt_0_4 = (_zz_cache_invld_gnt_0_3[7 : 4] | _zz_cache_invld_gnt_0_3[3 : 0]);
  assign cache_invld_gnt_0 = _zz_cache_invld_gnt_0_4[0];
  assign cache_invld_gnt_1 = _zz_cache_invld_gnt_0_4[1];
  assign cache_invld_gnt_2 = _zz_cache_invld_gnt_0_4[2];
  assign cache_invld_gnt_3 = _zz_cache_invld_gnt_0_4[3];
  assign _zz_cache_victim_gnt_0 = 4'b0001;
  assign _zz_cache_victim_gnt_0_1 = {cache_victim_3,{cache_victim_2,{cache_victim_1,cache_victim_0}}};
  assign _zz_cache_victim_gnt_0_2 = {_zz_cache_victim_gnt_0_1,_zz_cache_victim_gnt_0_1};
  assign _zz_cache_victim_gnt_0_3 = (_zz_cache_victim_gnt_0_2 & (~ _zz__zz_cache_victim_gnt_0_3));
  assign _zz_cache_victim_gnt_0_4 = (_zz_cache_victim_gnt_0_3[7 : 4] | _zz_cache_victim_gnt_0_3[3 : 0]);
  assign cache_victim_gnt_0 = _zz_cache_victim_gnt_0_4[0];
  assign cache_victim_gnt_1 = _zz_cache_victim_gnt_0_4[1];
  assign cache_victim_gnt_2 = _zz_cache_victim_gnt_0_4[2];
  assign cache_victim_gnt_3 = _zz_cache_victim_gnt_0_4[3];
  assign _zz_hit_id = (cache_hit_gnt_1 || cache_hit_gnt_3);
  assign _zz_hit_id_1 = (cache_hit_gnt_2 || cache_hit_gnt_3);
  assign hit_id = {_zz_hit_id_1,_zz_hit_id};
  assign _zz_invld_id = (cache_invld_gnt_1 || cache_invld_gnt_3);
  assign _zz_invld_id_1 = (cache_invld_gnt_2 || cache_invld_gnt_3);
  assign invld_id = {_zz_invld_id_1,_zz_invld_id};
  assign _zz_victim_id = (cache_victim_gnt_1 || cache_victim_gnt_3);
  assign _zz_victim_id_1 = (cache_victim_gnt_2 || cache_victim_gnt_3);
  assign victim_id = {_zz_victim_id_1,_zz_victim_id};
  assign evict_id = (is_diff ? invld_id : victim_id);
  assign _zz_1 = ({127'd0,1'b1} <<< cpu_set);
  assign _zz_2 = _zz_1[0];
  assign _zz_3 = _zz_1[1];
  assign _zz_4 = _zz_1[2];
  assign _zz_5 = _zz_1[3];
  assign _zz_6 = _zz_1[4];
  assign _zz_7 = _zz_1[5];
  assign _zz_8 = _zz_1[6];
  assign _zz_9 = _zz_1[7];
  assign _zz_10 = _zz_1[8];
  assign _zz_11 = _zz_1[9];
  assign _zz_12 = _zz_1[10];
  assign _zz_13 = _zz_1[11];
  assign _zz_14 = _zz_1[12];
  assign _zz_15 = _zz_1[13];
  assign _zz_16 = _zz_1[14];
  assign _zz_17 = _zz_1[15];
  assign _zz_18 = _zz_1[16];
  assign _zz_19 = _zz_1[17];
  assign _zz_20 = _zz_1[18];
  assign _zz_21 = _zz_1[19];
  assign _zz_22 = _zz_1[20];
  assign _zz_23 = _zz_1[21];
  assign _zz_24 = _zz_1[22];
  assign _zz_25 = _zz_1[23];
  assign _zz_26 = _zz_1[24];
  assign _zz_27 = _zz_1[25];
  assign _zz_28 = _zz_1[26];
  assign _zz_29 = _zz_1[27];
  assign _zz_30 = _zz_1[28];
  assign _zz_31 = _zz_1[29];
  assign _zz_32 = _zz_1[30];
  assign _zz_33 = _zz_1[31];
  assign _zz_34 = _zz_1[32];
  assign _zz_35 = _zz_1[33];
  assign _zz_36 = _zz_1[34];
  assign _zz_37 = _zz_1[35];
  assign _zz_38 = _zz_1[36];
  assign _zz_39 = _zz_1[37];
  assign _zz_40 = _zz_1[38];
  assign _zz_41 = _zz_1[39];
  assign _zz_42 = _zz_1[40];
  assign _zz_43 = _zz_1[41];
  assign _zz_44 = _zz_1[42];
  assign _zz_45 = _zz_1[43];
  assign _zz_46 = _zz_1[44];
  assign _zz_47 = _zz_1[45];
  assign _zz_48 = _zz_1[46];
  assign _zz_49 = _zz_1[47];
  assign _zz_50 = _zz_1[48];
  assign _zz_51 = _zz_1[49];
  assign _zz_52 = _zz_1[50];
  assign _zz_53 = _zz_1[51];
  assign _zz_54 = _zz_1[52];
  assign _zz_55 = _zz_1[53];
  assign _zz_56 = _zz_1[54];
  assign _zz_57 = _zz_1[55];
  assign _zz_58 = _zz_1[56];
  assign _zz_59 = _zz_1[57];
  assign _zz_60 = _zz_1[58];
  assign _zz_61 = _zz_1[59];
  assign _zz_62 = _zz_1[60];
  assign _zz_63 = _zz_1[61];
  assign _zz_64 = _zz_1[62];
  assign _zz_65 = _zz_1[63];
  assign _zz_66 = _zz_1[64];
  assign _zz_67 = _zz_1[65];
  assign _zz_68 = _zz_1[66];
  assign _zz_69 = _zz_1[67];
  assign _zz_70 = _zz_1[68];
  assign _zz_71 = _zz_1[69];
  assign _zz_72 = _zz_1[70];
  assign _zz_73 = _zz_1[71];
  assign _zz_74 = _zz_1[72];
  assign _zz_75 = _zz_1[73];
  assign _zz_76 = _zz_1[74];
  assign _zz_77 = _zz_1[75];
  assign _zz_78 = _zz_1[76];
  assign _zz_79 = _zz_1[77];
  assign _zz_80 = _zz_1[78];
  assign _zz_81 = _zz_1[79];
  assign _zz_82 = _zz_1[80];
  assign _zz_83 = _zz_1[81];
  assign _zz_84 = _zz_1[82];
  assign _zz_85 = _zz_1[83];
  assign _zz_86 = _zz_1[84];
  assign _zz_87 = _zz_1[85];
  assign _zz_88 = _zz_1[86];
  assign _zz_89 = _zz_1[87];
  assign _zz_90 = _zz_1[88];
  assign _zz_91 = _zz_1[89];
  assign _zz_92 = _zz_1[90];
  assign _zz_93 = _zz_1[91];
  assign _zz_94 = _zz_1[92];
  assign _zz_95 = _zz_1[93];
  assign _zz_96 = _zz_1[94];
  assign _zz_97 = _zz_1[95];
  assign _zz_98 = _zz_1[96];
  assign _zz_99 = _zz_1[97];
  assign _zz_100 = _zz_1[98];
  assign _zz_101 = _zz_1[99];
  assign _zz_102 = _zz_1[100];
  assign _zz_103 = _zz_1[101];
  assign _zz_104 = _zz_1[102];
  assign _zz_105 = _zz_1[103];
  assign _zz_106 = _zz_1[104];
  assign _zz_107 = _zz_1[105];
  assign _zz_108 = _zz_1[106];
  assign _zz_109 = _zz_1[107];
  assign _zz_110 = _zz_1[108];
  assign _zz_111 = _zz_1[109];
  assign _zz_112 = _zz_1[110];
  assign _zz_113 = _zz_1[111];
  assign _zz_114 = _zz_1[112];
  assign _zz_115 = _zz_1[113];
  assign _zz_116 = _zz_1[114];
  assign _zz_117 = _zz_1[115];
  assign _zz_118 = _zz_1[116];
  assign _zz_119 = _zz_1[117];
  assign _zz_120 = _zz_1[118];
  assign _zz_121 = _zz_1[119];
  assign _zz_122 = _zz_1[120];
  assign _zz_123 = _zz_1[121];
  assign _zz_124 = _zz_1[122];
  assign _zz_125 = _zz_1[123];
  assign _zz_126 = _zz_1[124];
  assign _zz_127 = _zz_1[125];
  assign _zz_128 = _zz_1[126];
  assign _zz_129 = _zz_1[127];
  assign cache_tag_0 = _zz_cache_tag_0;
  assign cache_hit_0 = ((cache_tag_0 == cpu_tag) && _zz_cache_hit_0);
  assign cache_mru_0 = _zz_cache_mru_0;
  assign _zz_130 = ({127'd0,1'b1} <<< cpu_set_d1);
  assign _zz_131 = _zz_130[0];
  assign _zz_132 = _zz_130[1];
  assign _zz_133 = _zz_130[2];
  assign _zz_134 = _zz_130[3];
  assign _zz_135 = _zz_130[4];
  assign _zz_136 = _zz_130[5];
  assign _zz_137 = _zz_130[6];
  assign _zz_138 = _zz_130[7];
  assign _zz_139 = _zz_130[8];
  assign _zz_140 = _zz_130[9];
  assign _zz_141 = _zz_130[10];
  assign _zz_142 = _zz_130[11];
  assign _zz_143 = _zz_130[12];
  assign _zz_144 = _zz_130[13];
  assign _zz_145 = _zz_130[14];
  assign _zz_146 = _zz_130[15];
  assign _zz_147 = _zz_130[16];
  assign _zz_148 = _zz_130[17];
  assign _zz_149 = _zz_130[18];
  assign _zz_150 = _zz_130[19];
  assign _zz_151 = _zz_130[20];
  assign _zz_152 = _zz_130[21];
  assign _zz_153 = _zz_130[22];
  assign _zz_154 = _zz_130[23];
  assign _zz_155 = _zz_130[24];
  assign _zz_156 = _zz_130[25];
  assign _zz_157 = _zz_130[26];
  assign _zz_158 = _zz_130[27];
  assign _zz_159 = _zz_130[28];
  assign _zz_160 = _zz_130[29];
  assign _zz_161 = _zz_130[30];
  assign _zz_162 = _zz_130[31];
  assign _zz_163 = _zz_130[32];
  assign _zz_164 = _zz_130[33];
  assign _zz_165 = _zz_130[34];
  assign _zz_166 = _zz_130[35];
  assign _zz_167 = _zz_130[36];
  assign _zz_168 = _zz_130[37];
  assign _zz_169 = _zz_130[38];
  assign _zz_170 = _zz_130[39];
  assign _zz_171 = _zz_130[40];
  assign _zz_172 = _zz_130[41];
  assign _zz_173 = _zz_130[42];
  assign _zz_174 = _zz_130[43];
  assign _zz_175 = _zz_130[44];
  assign _zz_176 = _zz_130[45];
  assign _zz_177 = _zz_130[46];
  assign _zz_178 = _zz_130[47];
  assign _zz_179 = _zz_130[48];
  assign _zz_180 = _zz_130[49];
  assign _zz_181 = _zz_130[50];
  assign _zz_182 = _zz_130[51];
  assign _zz_183 = _zz_130[52];
  assign _zz_184 = _zz_130[53];
  assign _zz_185 = _zz_130[54];
  assign _zz_186 = _zz_130[55];
  assign _zz_187 = _zz_130[56];
  assign _zz_188 = _zz_130[57];
  assign _zz_189 = _zz_130[58];
  assign _zz_190 = _zz_130[59];
  assign _zz_191 = _zz_130[60];
  assign _zz_192 = _zz_130[61];
  assign _zz_193 = _zz_130[62];
  assign _zz_194 = _zz_130[63];
  assign _zz_195 = _zz_130[64];
  assign _zz_196 = _zz_130[65];
  assign _zz_197 = _zz_130[66];
  assign _zz_198 = _zz_130[67];
  assign _zz_199 = _zz_130[68];
  assign _zz_200 = _zz_130[69];
  assign _zz_201 = _zz_130[70];
  assign _zz_202 = _zz_130[71];
  assign _zz_203 = _zz_130[72];
  assign _zz_204 = _zz_130[73];
  assign _zz_205 = _zz_130[74];
  assign _zz_206 = _zz_130[75];
  assign _zz_207 = _zz_130[76];
  assign _zz_208 = _zz_130[77];
  assign _zz_209 = _zz_130[78];
  assign _zz_210 = _zz_130[79];
  assign _zz_211 = _zz_130[80];
  assign _zz_212 = _zz_130[81];
  assign _zz_213 = _zz_130[82];
  assign _zz_214 = _zz_130[83];
  assign _zz_215 = _zz_130[84];
  assign _zz_216 = _zz_130[85];
  assign _zz_217 = _zz_130[86];
  assign _zz_218 = _zz_130[87];
  assign _zz_219 = _zz_130[88];
  assign _zz_220 = _zz_130[89];
  assign _zz_221 = _zz_130[90];
  assign _zz_222 = _zz_130[91];
  assign _zz_223 = _zz_130[92];
  assign _zz_224 = _zz_130[93];
  assign _zz_225 = _zz_130[94];
  assign _zz_226 = _zz_130[95];
  assign _zz_227 = _zz_130[96];
  assign _zz_228 = _zz_130[97];
  assign _zz_229 = _zz_130[98];
  assign _zz_230 = _zz_130[99];
  assign _zz_231 = _zz_130[100];
  assign _zz_232 = _zz_130[101];
  assign _zz_233 = _zz_130[102];
  assign _zz_234 = _zz_130[103];
  assign _zz_235 = _zz_130[104];
  assign _zz_236 = _zz_130[105];
  assign _zz_237 = _zz_130[106];
  assign _zz_238 = _zz_130[107];
  assign _zz_239 = _zz_130[108];
  assign _zz_240 = _zz_130[109];
  assign _zz_241 = _zz_130[110];
  assign _zz_242 = _zz_130[111];
  assign _zz_243 = _zz_130[112];
  assign _zz_244 = _zz_130[113];
  assign _zz_245 = _zz_130[114];
  assign _zz_246 = _zz_130[115];
  assign _zz_247 = _zz_130[116];
  assign _zz_248 = _zz_130[117];
  assign _zz_249 = _zz_130[118];
  assign _zz_250 = _zz_130[119];
  assign _zz_251 = _zz_130[120];
  assign _zz_252 = _zz_130[121];
  assign _zz_253 = _zz_130[122];
  assign _zz_254 = _zz_130[123];
  assign _zz_255 = _zz_130[124];
  assign _zz_256 = _zz_130[125];
  assign _zz_257 = _zz_130[126];
  assign _zz_258 = _zz_130[127];
  assign cache_invld_d1_0 = (! _zz_cache_invld_d1_0);
  assign cache_lru_d1_0 = (! _zz_cache_lru_d1_0);
  assign cache_victim_0 = (cache_invld_d1_0 && cache_lru_d1_0);
  assign sram_banks_data_0 = sram_0_ports_rsp_payload_data;
  assign sram_banks_valid_0 = sram_0_ports_rsp_valid;
  assign when_ICache_l174 = (is_hit && (2'b00 == hit_id));
  always @(*) begin
    if(when_ICache_l174) begin
      sram_0_ports_cmd_payload_addr = cpu_bank_addr;
    end else begin
      if(when_ICache_l181) begin
        sram_0_ports_cmd_payload_addr = cpu_bank_addr_d1;
      end else begin
        if(when_ICache_l188) begin
          sram_0_ports_cmd_payload_addr = next_level_bank_addr;
        end else begin
          sram_0_ports_cmd_payload_addr = 7'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l174) begin
      sram_0_ports_cmd_valid = 1'b1;
    end else begin
      if(when_ICache_l181) begin
        sram_0_ports_cmd_valid = 1'b1;
      end else begin
        if(when_ICache_l188) begin
          sram_0_ports_cmd_valid = 1'b1;
        end else begin
          sram_0_ports_cmd_valid = 1'b0;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l174) begin
      sram_0_ports_cmd_payload_wen = 16'h0;
    end else begin
      if(when_ICache_l181) begin
        sram_0_ports_cmd_payload_wen = 16'h0;
      end else begin
        if(when_ICache_l188) begin
          sram_0_ports_cmd_payload_wen = (_zz_sram_0_ports_cmd_payload_wen <<< _zz_sram_0_ports_cmd_payload_wen_1);
        end else begin
          sram_0_ports_cmd_payload_wen = 16'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l174) begin
      sram_0_ports_cmd_payload_wdata = 512'h0;
    end else begin
      if(when_ICache_l181) begin
        sram_0_ports_cmd_payload_wdata = 512'h0;
      end else begin
        if(when_ICache_l188) begin
          sram_0_ports_cmd_payload_wdata = ({448'h0,next_level_rsp_payload_data} <<< _zz_sram_0_ports_cmd_payload_wdata);
        end else begin
          sram_0_ports_cmd_payload_wdata = 512'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l174) begin
      sram_0_ports_cmd_payload_wstrb = 64'h0;
    end else begin
      if(when_ICache_l181) begin
        sram_0_ports_cmd_payload_wstrb = 64'h0;
      end else begin
        if(when_ICache_l188) begin
          sram_0_ports_cmd_payload_wstrb = ({56'h0,8'hff} <<< _zz_sram_0_ports_cmd_payload_wstrb);
        end else begin
          sram_0_ports_cmd_payload_wstrb = 64'h0;
        end
      end
    end
  end

  assign _zz_1549 = zz__zz_sram_0_ports_cmd_payload_wen(1'b0);
  always @(*) _zz_sram_0_ports_cmd_payload_wen = _zz_1549;
  assign when_ICache_l181 = (next_level_done && (2'b00 == evict_id_miss));
  assign when_ICache_l188 = (next_level_rsp_valid && (2'b00 == evict_id_miss));
  assign _zz_259 = ({127'd0,1'b1} <<< flush_cnt_value);
  assign _zz_260 = _zz_259[0];
  assign _zz_261 = _zz_259[1];
  assign _zz_262 = _zz_259[2];
  assign _zz_263 = _zz_259[3];
  assign _zz_264 = _zz_259[4];
  assign _zz_265 = _zz_259[5];
  assign _zz_266 = _zz_259[6];
  assign _zz_267 = _zz_259[7];
  assign _zz_268 = _zz_259[8];
  assign _zz_269 = _zz_259[9];
  assign _zz_270 = _zz_259[10];
  assign _zz_271 = _zz_259[11];
  assign _zz_272 = _zz_259[12];
  assign _zz_273 = _zz_259[13];
  assign _zz_274 = _zz_259[14];
  assign _zz_275 = _zz_259[15];
  assign _zz_276 = _zz_259[16];
  assign _zz_277 = _zz_259[17];
  assign _zz_278 = _zz_259[18];
  assign _zz_279 = _zz_259[19];
  assign _zz_280 = _zz_259[20];
  assign _zz_281 = _zz_259[21];
  assign _zz_282 = _zz_259[22];
  assign _zz_283 = _zz_259[23];
  assign _zz_284 = _zz_259[24];
  assign _zz_285 = _zz_259[25];
  assign _zz_286 = _zz_259[26];
  assign _zz_287 = _zz_259[27];
  assign _zz_288 = _zz_259[28];
  assign _zz_289 = _zz_259[29];
  assign _zz_290 = _zz_259[30];
  assign _zz_291 = _zz_259[31];
  assign _zz_292 = _zz_259[32];
  assign _zz_293 = _zz_259[33];
  assign _zz_294 = _zz_259[34];
  assign _zz_295 = _zz_259[35];
  assign _zz_296 = _zz_259[36];
  assign _zz_297 = _zz_259[37];
  assign _zz_298 = _zz_259[38];
  assign _zz_299 = _zz_259[39];
  assign _zz_300 = _zz_259[40];
  assign _zz_301 = _zz_259[41];
  assign _zz_302 = _zz_259[42];
  assign _zz_303 = _zz_259[43];
  assign _zz_304 = _zz_259[44];
  assign _zz_305 = _zz_259[45];
  assign _zz_306 = _zz_259[46];
  assign _zz_307 = _zz_259[47];
  assign _zz_308 = _zz_259[48];
  assign _zz_309 = _zz_259[49];
  assign _zz_310 = _zz_259[50];
  assign _zz_311 = _zz_259[51];
  assign _zz_312 = _zz_259[52];
  assign _zz_313 = _zz_259[53];
  assign _zz_314 = _zz_259[54];
  assign _zz_315 = _zz_259[55];
  assign _zz_316 = _zz_259[56];
  assign _zz_317 = _zz_259[57];
  assign _zz_318 = _zz_259[58];
  assign _zz_319 = _zz_259[59];
  assign _zz_320 = _zz_259[60];
  assign _zz_321 = _zz_259[61];
  assign _zz_322 = _zz_259[62];
  assign _zz_323 = _zz_259[63];
  assign _zz_324 = _zz_259[64];
  assign _zz_325 = _zz_259[65];
  assign _zz_326 = _zz_259[66];
  assign _zz_327 = _zz_259[67];
  assign _zz_328 = _zz_259[68];
  assign _zz_329 = _zz_259[69];
  assign _zz_330 = _zz_259[70];
  assign _zz_331 = _zz_259[71];
  assign _zz_332 = _zz_259[72];
  assign _zz_333 = _zz_259[73];
  assign _zz_334 = _zz_259[74];
  assign _zz_335 = _zz_259[75];
  assign _zz_336 = _zz_259[76];
  assign _zz_337 = _zz_259[77];
  assign _zz_338 = _zz_259[78];
  assign _zz_339 = _zz_259[79];
  assign _zz_340 = _zz_259[80];
  assign _zz_341 = _zz_259[81];
  assign _zz_342 = _zz_259[82];
  assign _zz_343 = _zz_259[83];
  assign _zz_344 = _zz_259[84];
  assign _zz_345 = _zz_259[85];
  assign _zz_346 = _zz_259[86];
  assign _zz_347 = _zz_259[87];
  assign _zz_348 = _zz_259[88];
  assign _zz_349 = _zz_259[89];
  assign _zz_350 = _zz_259[90];
  assign _zz_351 = _zz_259[91];
  assign _zz_352 = _zz_259[92];
  assign _zz_353 = _zz_259[93];
  assign _zz_354 = _zz_259[94];
  assign _zz_355 = _zz_259[95];
  assign _zz_356 = _zz_259[96];
  assign _zz_357 = _zz_259[97];
  assign _zz_358 = _zz_259[98];
  assign _zz_359 = _zz_259[99];
  assign _zz_360 = _zz_259[100];
  assign _zz_361 = _zz_259[101];
  assign _zz_362 = _zz_259[102];
  assign _zz_363 = _zz_259[103];
  assign _zz_364 = _zz_259[104];
  assign _zz_365 = _zz_259[105];
  assign _zz_366 = _zz_259[106];
  assign _zz_367 = _zz_259[107];
  assign _zz_368 = _zz_259[108];
  assign _zz_369 = _zz_259[109];
  assign _zz_370 = _zz_259[110];
  assign _zz_371 = _zz_259[111];
  assign _zz_372 = _zz_259[112];
  assign _zz_373 = _zz_259[113];
  assign _zz_374 = _zz_259[114];
  assign _zz_375 = _zz_259[115];
  assign _zz_376 = _zz_259[116];
  assign _zz_377 = _zz_259[117];
  assign _zz_378 = _zz_259[118];
  assign _zz_379 = _zz_259[119];
  assign _zz_380 = _zz_259[120];
  assign _zz_381 = _zz_259[121];
  assign _zz_382 = _zz_259[122];
  assign _zz_383 = _zz_259[123];
  assign _zz_384 = _zz_259[124];
  assign _zz_385 = _zz_259[125];
  assign _zz_386 = _zz_259[126];
  assign _zz_387 = _zz_259[127];
  assign when_ICache_l210 = (is_hit && mru_full);
  assign when_ICache_l217 = (is_hit && cache_hit_0);
  assign when_ICache_l220 = (next_level_done && (2'b00 == evict_id_miss));
  assign when_ICache_l225 = (next_level_done && (2'b00 == evict_id_miss));
  assign when_ICache_l230 = (flush || is_miss);
  assign when_ICache_l233 = (flush_done || next_level_done);
  assign _zz_388 = ({127'd0,1'b1} <<< cpu_set);
  assign _zz_389 = _zz_388[0];
  assign _zz_390 = _zz_388[1];
  assign _zz_391 = _zz_388[2];
  assign _zz_392 = _zz_388[3];
  assign _zz_393 = _zz_388[4];
  assign _zz_394 = _zz_388[5];
  assign _zz_395 = _zz_388[6];
  assign _zz_396 = _zz_388[7];
  assign _zz_397 = _zz_388[8];
  assign _zz_398 = _zz_388[9];
  assign _zz_399 = _zz_388[10];
  assign _zz_400 = _zz_388[11];
  assign _zz_401 = _zz_388[12];
  assign _zz_402 = _zz_388[13];
  assign _zz_403 = _zz_388[14];
  assign _zz_404 = _zz_388[15];
  assign _zz_405 = _zz_388[16];
  assign _zz_406 = _zz_388[17];
  assign _zz_407 = _zz_388[18];
  assign _zz_408 = _zz_388[19];
  assign _zz_409 = _zz_388[20];
  assign _zz_410 = _zz_388[21];
  assign _zz_411 = _zz_388[22];
  assign _zz_412 = _zz_388[23];
  assign _zz_413 = _zz_388[24];
  assign _zz_414 = _zz_388[25];
  assign _zz_415 = _zz_388[26];
  assign _zz_416 = _zz_388[27];
  assign _zz_417 = _zz_388[28];
  assign _zz_418 = _zz_388[29];
  assign _zz_419 = _zz_388[30];
  assign _zz_420 = _zz_388[31];
  assign _zz_421 = _zz_388[32];
  assign _zz_422 = _zz_388[33];
  assign _zz_423 = _zz_388[34];
  assign _zz_424 = _zz_388[35];
  assign _zz_425 = _zz_388[36];
  assign _zz_426 = _zz_388[37];
  assign _zz_427 = _zz_388[38];
  assign _zz_428 = _zz_388[39];
  assign _zz_429 = _zz_388[40];
  assign _zz_430 = _zz_388[41];
  assign _zz_431 = _zz_388[42];
  assign _zz_432 = _zz_388[43];
  assign _zz_433 = _zz_388[44];
  assign _zz_434 = _zz_388[45];
  assign _zz_435 = _zz_388[46];
  assign _zz_436 = _zz_388[47];
  assign _zz_437 = _zz_388[48];
  assign _zz_438 = _zz_388[49];
  assign _zz_439 = _zz_388[50];
  assign _zz_440 = _zz_388[51];
  assign _zz_441 = _zz_388[52];
  assign _zz_442 = _zz_388[53];
  assign _zz_443 = _zz_388[54];
  assign _zz_444 = _zz_388[55];
  assign _zz_445 = _zz_388[56];
  assign _zz_446 = _zz_388[57];
  assign _zz_447 = _zz_388[58];
  assign _zz_448 = _zz_388[59];
  assign _zz_449 = _zz_388[60];
  assign _zz_450 = _zz_388[61];
  assign _zz_451 = _zz_388[62];
  assign _zz_452 = _zz_388[63];
  assign _zz_453 = _zz_388[64];
  assign _zz_454 = _zz_388[65];
  assign _zz_455 = _zz_388[66];
  assign _zz_456 = _zz_388[67];
  assign _zz_457 = _zz_388[68];
  assign _zz_458 = _zz_388[69];
  assign _zz_459 = _zz_388[70];
  assign _zz_460 = _zz_388[71];
  assign _zz_461 = _zz_388[72];
  assign _zz_462 = _zz_388[73];
  assign _zz_463 = _zz_388[74];
  assign _zz_464 = _zz_388[75];
  assign _zz_465 = _zz_388[76];
  assign _zz_466 = _zz_388[77];
  assign _zz_467 = _zz_388[78];
  assign _zz_468 = _zz_388[79];
  assign _zz_469 = _zz_388[80];
  assign _zz_470 = _zz_388[81];
  assign _zz_471 = _zz_388[82];
  assign _zz_472 = _zz_388[83];
  assign _zz_473 = _zz_388[84];
  assign _zz_474 = _zz_388[85];
  assign _zz_475 = _zz_388[86];
  assign _zz_476 = _zz_388[87];
  assign _zz_477 = _zz_388[88];
  assign _zz_478 = _zz_388[89];
  assign _zz_479 = _zz_388[90];
  assign _zz_480 = _zz_388[91];
  assign _zz_481 = _zz_388[92];
  assign _zz_482 = _zz_388[93];
  assign _zz_483 = _zz_388[94];
  assign _zz_484 = _zz_388[95];
  assign _zz_485 = _zz_388[96];
  assign _zz_486 = _zz_388[97];
  assign _zz_487 = _zz_388[98];
  assign _zz_488 = _zz_388[99];
  assign _zz_489 = _zz_388[100];
  assign _zz_490 = _zz_388[101];
  assign _zz_491 = _zz_388[102];
  assign _zz_492 = _zz_388[103];
  assign _zz_493 = _zz_388[104];
  assign _zz_494 = _zz_388[105];
  assign _zz_495 = _zz_388[106];
  assign _zz_496 = _zz_388[107];
  assign _zz_497 = _zz_388[108];
  assign _zz_498 = _zz_388[109];
  assign _zz_499 = _zz_388[110];
  assign _zz_500 = _zz_388[111];
  assign _zz_501 = _zz_388[112];
  assign _zz_502 = _zz_388[113];
  assign _zz_503 = _zz_388[114];
  assign _zz_504 = _zz_388[115];
  assign _zz_505 = _zz_388[116];
  assign _zz_506 = _zz_388[117];
  assign _zz_507 = _zz_388[118];
  assign _zz_508 = _zz_388[119];
  assign _zz_509 = _zz_388[120];
  assign _zz_510 = _zz_388[121];
  assign _zz_511 = _zz_388[122];
  assign _zz_512 = _zz_388[123];
  assign _zz_513 = _zz_388[124];
  assign _zz_514 = _zz_388[125];
  assign _zz_515 = _zz_388[126];
  assign _zz_516 = _zz_388[127];
  assign cache_tag_1 = _zz_cache_tag_1;
  assign cache_hit_1 = ((cache_tag_1 == cpu_tag) && _zz_cache_hit_1);
  assign cache_mru_1 = _zz_cache_mru_1;
  assign _zz_517 = ({127'd0,1'b1} <<< cpu_set_d1);
  assign _zz_518 = _zz_517[0];
  assign _zz_519 = _zz_517[1];
  assign _zz_520 = _zz_517[2];
  assign _zz_521 = _zz_517[3];
  assign _zz_522 = _zz_517[4];
  assign _zz_523 = _zz_517[5];
  assign _zz_524 = _zz_517[6];
  assign _zz_525 = _zz_517[7];
  assign _zz_526 = _zz_517[8];
  assign _zz_527 = _zz_517[9];
  assign _zz_528 = _zz_517[10];
  assign _zz_529 = _zz_517[11];
  assign _zz_530 = _zz_517[12];
  assign _zz_531 = _zz_517[13];
  assign _zz_532 = _zz_517[14];
  assign _zz_533 = _zz_517[15];
  assign _zz_534 = _zz_517[16];
  assign _zz_535 = _zz_517[17];
  assign _zz_536 = _zz_517[18];
  assign _zz_537 = _zz_517[19];
  assign _zz_538 = _zz_517[20];
  assign _zz_539 = _zz_517[21];
  assign _zz_540 = _zz_517[22];
  assign _zz_541 = _zz_517[23];
  assign _zz_542 = _zz_517[24];
  assign _zz_543 = _zz_517[25];
  assign _zz_544 = _zz_517[26];
  assign _zz_545 = _zz_517[27];
  assign _zz_546 = _zz_517[28];
  assign _zz_547 = _zz_517[29];
  assign _zz_548 = _zz_517[30];
  assign _zz_549 = _zz_517[31];
  assign _zz_550 = _zz_517[32];
  assign _zz_551 = _zz_517[33];
  assign _zz_552 = _zz_517[34];
  assign _zz_553 = _zz_517[35];
  assign _zz_554 = _zz_517[36];
  assign _zz_555 = _zz_517[37];
  assign _zz_556 = _zz_517[38];
  assign _zz_557 = _zz_517[39];
  assign _zz_558 = _zz_517[40];
  assign _zz_559 = _zz_517[41];
  assign _zz_560 = _zz_517[42];
  assign _zz_561 = _zz_517[43];
  assign _zz_562 = _zz_517[44];
  assign _zz_563 = _zz_517[45];
  assign _zz_564 = _zz_517[46];
  assign _zz_565 = _zz_517[47];
  assign _zz_566 = _zz_517[48];
  assign _zz_567 = _zz_517[49];
  assign _zz_568 = _zz_517[50];
  assign _zz_569 = _zz_517[51];
  assign _zz_570 = _zz_517[52];
  assign _zz_571 = _zz_517[53];
  assign _zz_572 = _zz_517[54];
  assign _zz_573 = _zz_517[55];
  assign _zz_574 = _zz_517[56];
  assign _zz_575 = _zz_517[57];
  assign _zz_576 = _zz_517[58];
  assign _zz_577 = _zz_517[59];
  assign _zz_578 = _zz_517[60];
  assign _zz_579 = _zz_517[61];
  assign _zz_580 = _zz_517[62];
  assign _zz_581 = _zz_517[63];
  assign _zz_582 = _zz_517[64];
  assign _zz_583 = _zz_517[65];
  assign _zz_584 = _zz_517[66];
  assign _zz_585 = _zz_517[67];
  assign _zz_586 = _zz_517[68];
  assign _zz_587 = _zz_517[69];
  assign _zz_588 = _zz_517[70];
  assign _zz_589 = _zz_517[71];
  assign _zz_590 = _zz_517[72];
  assign _zz_591 = _zz_517[73];
  assign _zz_592 = _zz_517[74];
  assign _zz_593 = _zz_517[75];
  assign _zz_594 = _zz_517[76];
  assign _zz_595 = _zz_517[77];
  assign _zz_596 = _zz_517[78];
  assign _zz_597 = _zz_517[79];
  assign _zz_598 = _zz_517[80];
  assign _zz_599 = _zz_517[81];
  assign _zz_600 = _zz_517[82];
  assign _zz_601 = _zz_517[83];
  assign _zz_602 = _zz_517[84];
  assign _zz_603 = _zz_517[85];
  assign _zz_604 = _zz_517[86];
  assign _zz_605 = _zz_517[87];
  assign _zz_606 = _zz_517[88];
  assign _zz_607 = _zz_517[89];
  assign _zz_608 = _zz_517[90];
  assign _zz_609 = _zz_517[91];
  assign _zz_610 = _zz_517[92];
  assign _zz_611 = _zz_517[93];
  assign _zz_612 = _zz_517[94];
  assign _zz_613 = _zz_517[95];
  assign _zz_614 = _zz_517[96];
  assign _zz_615 = _zz_517[97];
  assign _zz_616 = _zz_517[98];
  assign _zz_617 = _zz_517[99];
  assign _zz_618 = _zz_517[100];
  assign _zz_619 = _zz_517[101];
  assign _zz_620 = _zz_517[102];
  assign _zz_621 = _zz_517[103];
  assign _zz_622 = _zz_517[104];
  assign _zz_623 = _zz_517[105];
  assign _zz_624 = _zz_517[106];
  assign _zz_625 = _zz_517[107];
  assign _zz_626 = _zz_517[108];
  assign _zz_627 = _zz_517[109];
  assign _zz_628 = _zz_517[110];
  assign _zz_629 = _zz_517[111];
  assign _zz_630 = _zz_517[112];
  assign _zz_631 = _zz_517[113];
  assign _zz_632 = _zz_517[114];
  assign _zz_633 = _zz_517[115];
  assign _zz_634 = _zz_517[116];
  assign _zz_635 = _zz_517[117];
  assign _zz_636 = _zz_517[118];
  assign _zz_637 = _zz_517[119];
  assign _zz_638 = _zz_517[120];
  assign _zz_639 = _zz_517[121];
  assign _zz_640 = _zz_517[122];
  assign _zz_641 = _zz_517[123];
  assign _zz_642 = _zz_517[124];
  assign _zz_643 = _zz_517[125];
  assign _zz_644 = _zz_517[126];
  assign _zz_645 = _zz_517[127];
  assign cache_invld_d1_1 = (! _zz_cache_invld_d1_1);
  assign cache_lru_d1_1 = (! _zz_cache_lru_d1_1);
  assign cache_victim_1 = (cache_invld_d1_1 && cache_lru_d1_1);
  assign sram_banks_data_1 = sram_1_ports_rsp_payload_data;
  assign sram_banks_valid_1 = sram_1_ports_rsp_valid;
  assign when_ICache_l174_1 = (is_hit && (2'b01 == hit_id));
  always @(*) begin
    if(when_ICache_l174_1) begin
      sram_1_ports_cmd_payload_addr = cpu_bank_addr;
    end else begin
      if(when_ICache_l181_1) begin
        sram_1_ports_cmd_payload_addr = cpu_bank_addr_d1;
      end else begin
        if(when_ICache_l188_1) begin
          sram_1_ports_cmd_payload_addr = next_level_bank_addr;
        end else begin
          sram_1_ports_cmd_payload_addr = 7'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l174_1) begin
      sram_1_ports_cmd_valid = 1'b1;
    end else begin
      if(when_ICache_l181_1) begin
        sram_1_ports_cmd_valid = 1'b1;
      end else begin
        if(when_ICache_l188_1) begin
          sram_1_ports_cmd_valid = 1'b1;
        end else begin
          sram_1_ports_cmd_valid = 1'b0;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l174_1) begin
      sram_1_ports_cmd_payload_wen = 16'h0;
    end else begin
      if(when_ICache_l181_1) begin
        sram_1_ports_cmd_payload_wen = 16'h0;
      end else begin
        if(when_ICache_l188_1) begin
          sram_1_ports_cmd_payload_wen = (_zz_sram_1_ports_cmd_payload_wen <<< _zz_sram_1_ports_cmd_payload_wen_1);
        end else begin
          sram_1_ports_cmd_payload_wen = 16'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l174_1) begin
      sram_1_ports_cmd_payload_wdata = 512'h0;
    end else begin
      if(when_ICache_l181_1) begin
        sram_1_ports_cmd_payload_wdata = 512'h0;
      end else begin
        if(when_ICache_l188_1) begin
          sram_1_ports_cmd_payload_wdata = ({448'h0,next_level_rsp_payload_data} <<< _zz_sram_1_ports_cmd_payload_wdata);
        end else begin
          sram_1_ports_cmd_payload_wdata = 512'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l174_1) begin
      sram_1_ports_cmd_payload_wstrb = 64'h0;
    end else begin
      if(when_ICache_l181_1) begin
        sram_1_ports_cmd_payload_wstrb = 64'h0;
      end else begin
        if(when_ICache_l188_1) begin
          sram_1_ports_cmd_payload_wstrb = ({56'h0,8'hff} <<< _zz_sram_1_ports_cmd_payload_wstrb);
        end else begin
          sram_1_ports_cmd_payload_wstrb = 64'h0;
        end
      end
    end
  end

  assign _zz_1550 = zz__zz_sram_1_ports_cmd_payload_wen(1'b0);
  always @(*) _zz_sram_1_ports_cmd_payload_wen = _zz_1550;
  assign when_ICache_l181_1 = (next_level_done && (2'b01 == evict_id_miss));
  assign when_ICache_l188_1 = (next_level_rsp_valid && (2'b01 == evict_id_miss));
  assign _zz_646 = ({127'd0,1'b1} <<< flush_cnt_value);
  assign _zz_647 = _zz_646[0];
  assign _zz_648 = _zz_646[1];
  assign _zz_649 = _zz_646[2];
  assign _zz_650 = _zz_646[3];
  assign _zz_651 = _zz_646[4];
  assign _zz_652 = _zz_646[5];
  assign _zz_653 = _zz_646[6];
  assign _zz_654 = _zz_646[7];
  assign _zz_655 = _zz_646[8];
  assign _zz_656 = _zz_646[9];
  assign _zz_657 = _zz_646[10];
  assign _zz_658 = _zz_646[11];
  assign _zz_659 = _zz_646[12];
  assign _zz_660 = _zz_646[13];
  assign _zz_661 = _zz_646[14];
  assign _zz_662 = _zz_646[15];
  assign _zz_663 = _zz_646[16];
  assign _zz_664 = _zz_646[17];
  assign _zz_665 = _zz_646[18];
  assign _zz_666 = _zz_646[19];
  assign _zz_667 = _zz_646[20];
  assign _zz_668 = _zz_646[21];
  assign _zz_669 = _zz_646[22];
  assign _zz_670 = _zz_646[23];
  assign _zz_671 = _zz_646[24];
  assign _zz_672 = _zz_646[25];
  assign _zz_673 = _zz_646[26];
  assign _zz_674 = _zz_646[27];
  assign _zz_675 = _zz_646[28];
  assign _zz_676 = _zz_646[29];
  assign _zz_677 = _zz_646[30];
  assign _zz_678 = _zz_646[31];
  assign _zz_679 = _zz_646[32];
  assign _zz_680 = _zz_646[33];
  assign _zz_681 = _zz_646[34];
  assign _zz_682 = _zz_646[35];
  assign _zz_683 = _zz_646[36];
  assign _zz_684 = _zz_646[37];
  assign _zz_685 = _zz_646[38];
  assign _zz_686 = _zz_646[39];
  assign _zz_687 = _zz_646[40];
  assign _zz_688 = _zz_646[41];
  assign _zz_689 = _zz_646[42];
  assign _zz_690 = _zz_646[43];
  assign _zz_691 = _zz_646[44];
  assign _zz_692 = _zz_646[45];
  assign _zz_693 = _zz_646[46];
  assign _zz_694 = _zz_646[47];
  assign _zz_695 = _zz_646[48];
  assign _zz_696 = _zz_646[49];
  assign _zz_697 = _zz_646[50];
  assign _zz_698 = _zz_646[51];
  assign _zz_699 = _zz_646[52];
  assign _zz_700 = _zz_646[53];
  assign _zz_701 = _zz_646[54];
  assign _zz_702 = _zz_646[55];
  assign _zz_703 = _zz_646[56];
  assign _zz_704 = _zz_646[57];
  assign _zz_705 = _zz_646[58];
  assign _zz_706 = _zz_646[59];
  assign _zz_707 = _zz_646[60];
  assign _zz_708 = _zz_646[61];
  assign _zz_709 = _zz_646[62];
  assign _zz_710 = _zz_646[63];
  assign _zz_711 = _zz_646[64];
  assign _zz_712 = _zz_646[65];
  assign _zz_713 = _zz_646[66];
  assign _zz_714 = _zz_646[67];
  assign _zz_715 = _zz_646[68];
  assign _zz_716 = _zz_646[69];
  assign _zz_717 = _zz_646[70];
  assign _zz_718 = _zz_646[71];
  assign _zz_719 = _zz_646[72];
  assign _zz_720 = _zz_646[73];
  assign _zz_721 = _zz_646[74];
  assign _zz_722 = _zz_646[75];
  assign _zz_723 = _zz_646[76];
  assign _zz_724 = _zz_646[77];
  assign _zz_725 = _zz_646[78];
  assign _zz_726 = _zz_646[79];
  assign _zz_727 = _zz_646[80];
  assign _zz_728 = _zz_646[81];
  assign _zz_729 = _zz_646[82];
  assign _zz_730 = _zz_646[83];
  assign _zz_731 = _zz_646[84];
  assign _zz_732 = _zz_646[85];
  assign _zz_733 = _zz_646[86];
  assign _zz_734 = _zz_646[87];
  assign _zz_735 = _zz_646[88];
  assign _zz_736 = _zz_646[89];
  assign _zz_737 = _zz_646[90];
  assign _zz_738 = _zz_646[91];
  assign _zz_739 = _zz_646[92];
  assign _zz_740 = _zz_646[93];
  assign _zz_741 = _zz_646[94];
  assign _zz_742 = _zz_646[95];
  assign _zz_743 = _zz_646[96];
  assign _zz_744 = _zz_646[97];
  assign _zz_745 = _zz_646[98];
  assign _zz_746 = _zz_646[99];
  assign _zz_747 = _zz_646[100];
  assign _zz_748 = _zz_646[101];
  assign _zz_749 = _zz_646[102];
  assign _zz_750 = _zz_646[103];
  assign _zz_751 = _zz_646[104];
  assign _zz_752 = _zz_646[105];
  assign _zz_753 = _zz_646[106];
  assign _zz_754 = _zz_646[107];
  assign _zz_755 = _zz_646[108];
  assign _zz_756 = _zz_646[109];
  assign _zz_757 = _zz_646[110];
  assign _zz_758 = _zz_646[111];
  assign _zz_759 = _zz_646[112];
  assign _zz_760 = _zz_646[113];
  assign _zz_761 = _zz_646[114];
  assign _zz_762 = _zz_646[115];
  assign _zz_763 = _zz_646[116];
  assign _zz_764 = _zz_646[117];
  assign _zz_765 = _zz_646[118];
  assign _zz_766 = _zz_646[119];
  assign _zz_767 = _zz_646[120];
  assign _zz_768 = _zz_646[121];
  assign _zz_769 = _zz_646[122];
  assign _zz_770 = _zz_646[123];
  assign _zz_771 = _zz_646[124];
  assign _zz_772 = _zz_646[125];
  assign _zz_773 = _zz_646[126];
  assign _zz_774 = _zz_646[127];
  assign when_ICache_l210_1 = (is_hit && mru_full);
  assign when_ICache_l217_1 = (is_hit && cache_hit_1);
  assign when_ICache_l220_1 = (next_level_done && (2'b01 == evict_id_miss));
  assign when_ICache_l225_1 = (next_level_done && (2'b01 == evict_id_miss));
  assign when_ICache_l230_1 = (flush || is_miss);
  assign when_ICache_l233_1 = (flush_done || next_level_done);
  assign _zz_775 = ({127'd0,1'b1} <<< cpu_set);
  assign _zz_776 = _zz_775[0];
  assign _zz_777 = _zz_775[1];
  assign _zz_778 = _zz_775[2];
  assign _zz_779 = _zz_775[3];
  assign _zz_780 = _zz_775[4];
  assign _zz_781 = _zz_775[5];
  assign _zz_782 = _zz_775[6];
  assign _zz_783 = _zz_775[7];
  assign _zz_784 = _zz_775[8];
  assign _zz_785 = _zz_775[9];
  assign _zz_786 = _zz_775[10];
  assign _zz_787 = _zz_775[11];
  assign _zz_788 = _zz_775[12];
  assign _zz_789 = _zz_775[13];
  assign _zz_790 = _zz_775[14];
  assign _zz_791 = _zz_775[15];
  assign _zz_792 = _zz_775[16];
  assign _zz_793 = _zz_775[17];
  assign _zz_794 = _zz_775[18];
  assign _zz_795 = _zz_775[19];
  assign _zz_796 = _zz_775[20];
  assign _zz_797 = _zz_775[21];
  assign _zz_798 = _zz_775[22];
  assign _zz_799 = _zz_775[23];
  assign _zz_800 = _zz_775[24];
  assign _zz_801 = _zz_775[25];
  assign _zz_802 = _zz_775[26];
  assign _zz_803 = _zz_775[27];
  assign _zz_804 = _zz_775[28];
  assign _zz_805 = _zz_775[29];
  assign _zz_806 = _zz_775[30];
  assign _zz_807 = _zz_775[31];
  assign _zz_808 = _zz_775[32];
  assign _zz_809 = _zz_775[33];
  assign _zz_810 = _zz_775[34];
  assign _zz_811 = _zz_775[35];
  assign _zz_812 = _zz_775[36];
  assign _zz_813 = _zz_775[37];
  assign _zz_814 = _zz_775[38];
  assign _zz_815 = _zz_775[39];
  assign _zz_816 = _zz_775[40];
  assign _zz_817 = _zz_775[41];
  assign _zz_818 = _zz_775[42];
  assign _zz_819 = _zz_775[43];
  assign _zz_820 = _zz_775[44];
  assign _zz_821 = _zz_775[45];
  assign _zz_822 = _zz_775[46];
  assign _zz_823 = _zz_775[47];
  assign _zz_824 = _zz_775[48];
  assign _zz_825 = _zz_775[49];
  assign _zz_826 = _zz_775[50];
  assign _zz_827 = _zz_775[51];
  assign _zz_828 = _zz_775[52];
  assign _zz_829 = _zz_775[53];
  assign _zz_830 = _zz_775[54];
  assign _zz_831 = _zz_775[55];
  assign _zz_832 = _zz_775[56];
  assign _zz_833 = _zz_775[57];
  assign _zz_834 = _zz_775[58];
  assign _zz_835 = _zz_775[59];
  assign _zz_836 = _zz_775[60];
  assign _zz_837 = _zz_775[61];
  assign _zz_838 = _zz_775[62];
  assign _zz_839 = _zz_775[63];
  assign _zz_840 = _zz_775[64];
  assign _zz_841 = _zz_775[65];
  assign _zz_842 = _zz_775[66];
  assign _zz_843 = _zz_775[67];
  assign _zz_844 = _zz_775[68];
  assign _zz_845 = _zz_775[69];
  assign _zz_846 = _zz_775[70];
  assign _zz_847 = _zz_775[71];
  assign _zz_848 = _zz_775[72];
  assign _zz_849 = _zz_775[73];
  assign _zz_850 = _zz_775[74];
  assign _zz_851 = _zz_775[75];
  assign _zz_852 = _zz_775[76];
  assign _zz_853 = _zz_775[77];
  assign _zz_854 = _zz_775[78];
  assign _zz_855 = _zz_775[79];
  assign _zz_856 = _zz_775[80];
  assign _zz_857 = _zz_775[81];
  assign _zz_858 = _zz_775[82];
  assign _zz_859 = _zz_775[83];
  assign _zz_860 = _zz_775[84];
  assign _zz_861 = _zz_775[85];
  assign _zz_862 = _zz_775[86];
  assign _zz_863 = _zz_775[87];
  assign _zz_864 = _zz_775[88];
  assign _zz_865 = _zz_775[89];
  assign _zz_866 = _zz_775[90];
  assign _zz_867 = _zz_775[91];
  assign _zz_868 = _zz_775[92];
  assign _zz_869 = _zz_775[93];
  assign _zz_870 = _zz_775[94];
  assign _zz_871 = _zz_775[95];
  assign _zz_872 = _zz_775[96];
  assign _zz_873 = _zz_775[97];
  assign _zz_874 = _zz_775[98];
  assign _zz_875 = _zz_775[99];
  assign _zz_876 = _zz_775[100];
  assign _zz_877 = _zz_775[101];
  assign _zz_878 = _zz_775[102];
  assign _zz_879 = _zz_775[103];
  assign _zz_880 = _zz_775[104];
  assign _zz_881 = _zz_775[105];
  assign _zz_882 = _zz_775[106];
  assign _zz_883 = _zz_775[107];
  assign _zz_884 = _zz_775[108];
  assign _zz_885 = _zz_775[109];
  assign _zz_886 = _zz_775[110];
  assign _zz_887 = _zz_775[111];
  assign _zz_888 = _zz_775[112];
  assign _zz_889 = _zz_775[113];
  assign _zz_890 = _zz_775[114];
  assign _zz_891 = _zz_775[115];
  assign _zz_892 = _zz_775[116];
  assign _zz_893 = _zz_775[117];
  assign _zz_894 = _zz_775[118];
  assign _zz_895 = _zz_775[119];
  assign _zz_896 = _zz_775[120];
  assign _zz_897 = _zz_775[121];
  assign _zz_898 = _zz_775[122];
  assign _zz_899 = _zz_775[123];
  assign _zz_900 = _zz_775[124];
  assign _zz_901 = _zz_775[125];
  assign _zz_902 = _zz_775[126];
  assign _zz_903 = _zz_775[127];
  assign cache_tag_2 = _zz_cache_tag_2;
  assign cache_hit_2 = ((cache_tag_2 == cpu_tag) && _zz_cache_hit_2);
  assign cache_mru_2 = _zz_cache_mru_2;
  assign _zz_904 = ({127'd0,1'b1} <<< cpu_set_d1);
  assign _zz_905 = _zz_904[0];
  assign _zz_906 = _zz_904[1];
  assign _zz_907 = _zz_904[2];
  assign _zz_908 = _zz_904[3];
  assign _zz_909 = _zz_904[4];
  assign _zz_910 = _zz_904[5];
  assign _zz_911 = _zz_904[6];
  assign _zz_912 = _zz_904[7];
  assign _zz_913 = _zz_904[8];
  assign _zz_914 = _zz_904[9];
  assign _zz_915 = _zz_904[10];
  assign _zz_916 = _zz_904[11];
  assign _zz_917 = _zz_904[12];
  assign _zz_918 = _zz_904[13];
  assign _zz_919 = _zz_904[14];
  assign _zz_920 = _zz_904[15];
  assign _zz_921 = _zz_904[16];
  assign _zz_922 = _zz_904[17];
  assign _zz_923 = _zz_904[18];
  assign _zz_924 = _zz_904[19];
  assign _zz_925 = _zz_904[20];
  assign _zz_926 = _zz_904[21];
  assign _zz_927 = _zz_904[22];
  assign _zz_928 = _zz_904[23];
  assign _zz_929 = _zz_904[24];
  assign _zz_930 = _zz_904[25];
  assign _zz_931 = _zz_904[26];
  assign _zz_932 = _zz_904[27];
  assign _zz_933 = _zz_904[28];
  assign _zz_934 = _zz_904[29];
  assign _zz_935 = _zz_904[30];
  assign _zz_936 = _zz_904[31];
  assign _zz_937 = _zz_904[32];
  assign _zz_938 = _zz_904[33];
  assign _zz_939 = _zz_904[34];
  assign _zz_940 = _zz_904[35];
  assign _zz_941 = _zz_904[36];
  assign _zz_942 = _zz_904[37];
  assign _zz_943 = _zz_904[38];
  assign _zz_944 = _zz_904[39];
  assign _zz_945 = _zz_904[40];
  assign _zz_946 = _zz_904[41];
  assign _zz_947 = _zz_904[42];
  assign _zz_948 = _zz_904[43];
  assign _zz_949 = _zz_904[44];
  assign _zz_950 = _zz_904[45];
  assign _zz_951 = _zz_904[46];
  assign _zz_952 = _zz_904[47];
  assign _zz_953 = _zz_904[48];
  assign _zz_954 = _zz_904[49];
  assign _zz_955 = _zz_904[50];
  assign _zz_956 = _zz_904[51];
  assign _zz_957 = _zz_904[52];
  assign _zz_958 = _zz_904[53];
  assign _zz_959 = _zz_904[54];
  assign _zz_960 = _zz_904[55];
  assign _zz_961 = _zz_904[56];
  assign _zz_962 = _zz_904[57];
  assign _zz_963 = _zz_904[58];
  assign _zz_964 = _zz_904[59];
  assign _zz_965 = _zz_904[60];
  assign _zz_966 = _zz_904[61];
  assign _zz_967 = _zz_904[62];
  assign _zz_968 = _zz_904[63];
  assign _zz_969 = _zz_904[64];
  assign _zz_970 = _zz_904[65];
  assign _zz_971 = _zz_904[66];
  assign _zz_972 = _zz_904[67];
  assign _zz_973 = _zz_904[68];
  assign _zz_974 = _zz_904[69];
  assign _zz_975 = _zz_904[70];
  assign _zz_976 = _zz_904[71];
  assign _zz_977 = _zz_904[72];
  assign _zz_978 = _zz_904[73];
  assign _zz_979 = _zz_904[74];
  assign _zz_980 = _zz_904[75];
  assign _zz_981 = _zz_904[76];
  assign _zz_982 = _zz_904[77];
  assign _zz_983 = _zz_904[78];
  assign _zz_984 = _zz_904[79];
  assign _zz_985 = _zz_904[80];
  assign _zz_986 = _zz_904[81];
  assign _zz_987 = _zz_904[82];
  assign _zz_988 = _zz_904[83];
  assign _zz_989 = _zz_904[84];
  assign _zz_990 = _zz_904[85];
  assign _zz_991 = _zz_904[86];
  assign _zz_992 = _zz_904[87];
  assign _zz_993 = _zz_904[88];
  assign _zz_994 = _zz_904[89];
  assign _zz_995 = _zz_904[90];
  assign _zz_996 = _zz_904[91];
  assign _zz_997 = _zz_904[92];
  assign _zz_998 = _zz_904[93];
  assign _zz_999 = _zz_904[94];
  assign _zz_1000 = _zz_904[95];
  assign _zz_1001 = _zz_904[96];
  assign _zz_1002 = _zz_904[97];
  assign _zz_1003 = _zz_904[98];
  assign _zz_1004 = _zz_904[99];
  assign _zz_1005 = _zz_904[100];
  assign _zz_1006 = _zz_904[101];
  assign _zz_1007 = _zz_904[102];
  assign _zz_1008 = _zz_904[103];
  assign _zz_1009 = _zz_904[104];
  assign _zz_1010 = _zz_904[105];
  assign _zz_1011 = _zz_904[106];
  assign _zz_1012 = _zz_904[107];
  assign _zz_1013 = _zz_904[108];
  assign _zz_1014 = _zz_904[109];
  assign _zz_1015 = _zz_904[110];
  assign _zz_1016 = _zz_904[111];
  assign _zz_1017 = _zz_904[112];
  assign _zz_1018 = _zz_904[113];
  assign _zz_1019 = _zz_904[114];
  assign _zz_1020 = _zz_904[115];
  assign _zz_1021 = _zz_904[116];
  assign _zz_1022 = _zz_904[117];
  assign _zz_1023 = _zz_904[118];
  assign _zz_1024 = _zz_904[119];
  assign _zz_1025 = _zz_904[120];
  assign _zz_1026 = _zz_904[121];
  assign _zz_1027 = _zz_904[122];
  assign _zz_1028 = _zz_904[123];
  assign _zz_1029 = _zz_904[124];
  assign _zz_1030 = _zz_904[125];
  assign _zz_1031 = _zz_904[126];
  assign _zz_1032 = _zz_904[127];
  assign cache_invld_d1_2 = (! _zz_cache_invld_d1_2);
  assign cache_lru_d1_2 = (! _zz_cache_lru_d1_2);
  assign cache_victim_2 = (cache_invld_d1_2 && cache_lru_d1_2);
  assign sram_banks_data_2 = sram_2_ports_rsp_payload_data;
  assign sram_banks_valid_2 = sram_2_ports_rsp_valid;
  assign when_ICache_l174_2 = (is_hit && (2'b10 == hit_id));
  always @(*) begin
    if(when_ICache_l174_2) begin
      sram_2_ports_cmd_payload_addr = cpu_bank_addr;
    end else begin
      if(when_ICache_l181_2) begin
        sram_2_ports_cmd_payload_addr = cpu_bank_addr_d1;
      end else begin
        if(when_ICache_l188_2) begin
          sram_2_ports_cmd_payload_addr = next_level_bank_addr;
        end else begin
          sram_2_ports_cmd_payload_addr = 7'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l174_2) begin
      sram_2_ports_cmd_valid = 1'b1;
    end else begin
      if(when_ICache_l181_2) begin
        sram_2_ports_cmd_valid = 1'b1;
      end else begin
        if(when_ICache_l188_2) begin
          sram_2_ports_cmd_valid = 1'b1;
        end else begin
          sram_2_ports_cmd_valid = 1'b0;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l174_2) begin
      sram_2_ports_cmd_payload_wen = 16'h0;
    end else begin
      if(when_ICache_l181_2) begin
        sram_2_ports_cmd_payload_wen = 16'h0;
      end else begin
        if(when_ICache_l188_2) begin
          sram_2_ports_cmd_payload_wen = (_zz_sram_2_ports_cmd_payload_wen <<< _zz_sram_2_ports_cmd_payload_wen_1);
        end else begin
          sram_2_ports_cmd_payload_wen = 16'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l174_2) begin
      sram_2_ports_cmd_payload_wdata = 512'h0;
    end else begin
      if(when_ICache_l181_2) begin
        sram_2_ports_cmd_payload_wdata = 512'h0;
      end else begin
        if(when_ICache_l188_2) begin
          sram_2_ports_cmd_payload_wdata = ({448'h0,next_level_rsp_payload_data} <<< _zz_sram_2_ports_cmd_payload_wdata);
        end else begin
          sram_2_ports_cmd_payload_wdata = 512'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l174_2) begin
      sram_2_ports_cmd_payload_wstrb = 64'h0;
    end else begin
      if(when_ICache_l181_2) begin
        sram_2_ports_cmd_payload_wstrb = 64'h0;
      end else begin
        if(when_ICache_l188_2) begin
          sram_2_ports_cmd_payload_wstrb = ({56'h0,8'hff} <<< _zz_sram_2_ports_cmd_payload_wstrb);
        end else begin
          sram_2_ports_cmd_payload_wstrb = 64'h0;
        end
      end
    end
  end

  assign _zz_1551 = zz__zz_sram_2_ports_cmd_payload_wen(1'b0);
  always @(*) _zz_sram_2_ports_cmd_payload_wen = _zz_1551;
  assign when_ICache_l181_2 = (next_level_done && (2'b10 == evict_id_miss));
  assign when_ICache_l188_2 = (next_level_rsp_valid && (2'b10 == evict_id_miss));
  assign _zz_1033 = ({127'd0,1'b1} <<< flush_cnt_value);
  assign _zz_1034 = _zz_1033[0];
  assign _zz_1035 = _zz_1033[1];
  assign _zz_1036 = _zz_1033[2];
  assign _zz_1037 = _zz_1033[3];
  assign _zz_1038 = _zz_1033[4];
  assign _zz_1039 = _zz_1033[5];
  assign _zz_1040 = _zz_1033[6];
  assign _zz_1041 = _zz_1033[7];
  assign _zz_1042 = _zz_1033[8];
  assign _zz_1043 = _zz_1033[9];
  assign _zz_1044 = _zz_1033[10];
  assign _zz_1045 = _zz_1033[11];
  assign _zz_1046 = _zz_1033[12];
  assign _zz_1047 = _zz_1033[13];
  assign _zz_1048 = _zz_1033[14];
  assign _zz_1049 = _zz_1033[15];
  assign _zz_1050 = _zz_1033[16];
  assign _zz_1051 = _zz_1033[17];
  assign _zz_1052 = _zz_1033[18];
  assign _zz_1053 = _zz_1033[19];
  assign _zz_1054 = _zz_1033[20];
  assign _zz_1055 = _zz_1033[21];
  assign _zz_1056 = _zz_1033[22];
  assign _zz_1057 = _zz_1033[23];
  assign _zz_1058 = _zz_1033[24];
  assign _zz_1059 = _zz_1033[25];
  assign _zz_1060 = _zz_1033[26];
  assign _zz_1061 = _zz_1033[27];
  assign _zz_1062 = _zz_1033[28];
  assign _zz_1063 = _zz_1033[29];
  assign _zz_1064 = _zz_1033[30];
  assign _zz_1065 = _zz_1033[31];
  assign _zz_1066 = _zz_1033[32];
  assign _zz_1067 = _zz_1033[33];
  assign _zz_1068 = _zz_1033[34];
  assign _zz_1069 = _zz_1033[35];
  assign _zz_1070 = _zz_1033[36];
  assign _zz_1071 = _zz_1033[37];
  assign _zz_1072 = _zz_1033[38];
  assign _zz_1073 = _zz_1033[39];
  assign _zz_1074 = _zz_1033[40];
  assign _zz_1075 = _zz_1033[41];
  assign _zz_1076 = _zz_1033[42];
  assign _zz_1077 = _zz_1033[43];
  assign _zz_1078 = _zz_1033[44];
  assign _zz_1079 = _zz_1033[45];
  assign _zz_1080 = _zz_1033[46];
  assign _zz_1081 = _zz_1033[47];
  assign _zz_1082 = _zz_1033[48];
  assign _zz_1083 = _zz_1033[49];
  assign _zz_1084 = _zz_1033[50];
  assign _zz_1085 = _zz_1033[51];
  assign _zz_1086 = _zz_1033[52];
  assign _zz_1087 = _zz_1033[53];
  assign _zz_1088 = _zz_1033[54];
  assign _zz_1089 = _zz_1033[55];
  assign _zz_1090 = _zz_1033[56];
  assign _zz_1091 = _zz_1033[57];
  assign _zz_1092 = _zz_1033[58];
  assign _zz_1093 = _zz_1033[59];
  assign _zz_1094 = _zz_1033[60];
  assign _zz_1095 = _zz_1033[61];
  assign _zz_1096 = _zz_1033[62];
  assign _zz_1097 = _zz_1033[63];
  assign _zz_1098 = _zz_1033[64];
  assign _zz_1099 = _zz_1033[65];
  assign _zz_1100 = _zz_1033[66];
  assign _zz_1101 = _zz_1033[67];
  assign _zz_1102 = _zz_1033[68];
  assign _zz_1103 = _zz_1033[69];
  assign _zz_1104 = _zz_1033[70];
  assign _zz_1105 = _zz_1033[71];
  assign _zz_1106 = _zz_1033[72];
  assign _zz_1107 = _zz_1033[73];
  assign _zz_1108 = _zz_1033[74];
  assign _zz_1109 = _zz_1033[75];
  assign _zz_1110 = _zz_1033[76];
  assign _zz_1111 = _zz_1033[77];
  assign _zz_1112 = _zz_1033[78];
  assign _zz_1113 = _zz_1033[79];
  assign _zz_1114 = _zz_1033[80];
  assign _zz_1115 = _zz_1033[81];
  assign _zz_1116 = _zz_1033[82];
  assign _zz_1117 = _zz_1033[83];
  assign _zz_1118 = _zz_1033[84];
  assign _zz_1119 = _zz_1033[85];
  assign _zz_1120 = _zz_1033[86];
  assign _zz_1121 = _zz_1033[87];
  assign _zz_1122 = _zz_1033[88];
  assign _zz_1123 = _zz_1033[89];
  assign _zz_1124 = _zz_1033[90];
  assign _zz_1125 = _zz_1033[91];
  assign _zz_1126 = _zz_1033[92];
  assign _zz_1127 = _zz_1033[93];
  assign _zz_1128 = _zz_1033[94];
  assign _zz_1129 = _zz_1033[95];
  assign _zz_1130 = _zz_1033[96];
  assign _zz_1131 = _zz_1033[97];
  assign _zz_1132 = _zz_1033[98];
  assign _zz_1133 = _zz_1033[99];
  assign _zz_1134 = _zz_1033[100];
  assign _zz_1135 = _zz_1033[101];
  assign _zz_1136 = _zz_1033[102];
  assign _zz_1137 = _zz_1033[103];
  assign _zz_1138 = _zz_1033[104];
  assign _zz_1139 = _zz_1033[105];
  assign _zz_1140 = _zz_1033[106];
  assign _zz_1141 = _zz_1033[107];
  assign _zz_1142 = _zz_1033[108];
  assign _zz_1143 = _zz_1033[109];
  assign _zz_1144 = _zz_1033[110];
  assign _zz_1145 = _zz_1033[111];
  assign _zz_1146 = _zz_1033[112];
  assign _zz_1147 = _zz_1033[113];
  assign _zz_1148 = _zz_1033[114];
  assign _zz_1149 = _zz_1033[115];
  assign _zz_1150 = _zz_1033[116];
  assign _zz_1151 = _zz_1033[117];
  assign _zz_1152 = _zz_1033[118];
  assign _zz_1153 = _zz_1033[119];
  assign _zz_1154 = _zz_1033[120];
  assign _zz_1155 = _zz_1033[121];
  assign _zz_1156 = _zz_1033[122];
  assign _zz_1157 = _zz_1033[123];
  assign _zz_1158 = _zz_1033[124];
  assign _zz_1159 = _zz_1033[125];
  assign _zz_1160 = _zz_1033[126];
  assign _zz_1161 = _zz_1033[127];
  assign when_ICache_l210_2 = (is_hit && mru_full);
  assign when_ICache_l217_2 = (is_hit && cache_hit_2);
  assign when_ICache_l220_2 = (next_level_done && (2'b10 == evict_id_miss));
  assign when_ICache_l225_2 = (next_level_done && (2'b10 == evict_id_miss));
  assign when_ICache_l230_2 = (flush || is_miss);
  assign when_ICache_l233_2 = (flush_done || next_level_done);
  assign _zz_1162 = ({127'd0,1'b1} <<< cpu_set);
  assign _zz_1163 = _zz_1162[0];
  assign _zz_1164 = _zz_1162[1];
  assign _zz_1165 = _zz_1162[2];
  assign _zz_1166 = _zz_1162[3];
  assign _zz_1167 = _zz_1162[4];
  assign _zz_1168 = _zz_1162[5];
  assign _zz_1169 = _zz_1162[6];
  assign _zz_1170 = _zz_1162[7];
  assign _zz_1171 = _zz_1162[8];
  assign _zz_1172 = _zz_1162[9];
  assign _zz_1173 = _zz_1162[10];
  assign _zz_1174 = _zz_1162[11];
  assign _zz_1175 = _zz_1162[12];
  assign _zz_1176 = _zz_1162[13];
  assign _zz_1177 = _zz_1162[14];
  assign _zz_1178 = _zz_1162[15];
  assign _zz_1179 = _zz_1162[16];
  assign _zz_1180 = _zz_1162[17];
  assign _zz_1181 = _zz_1162[18];
  assign _zz_1182 = _zz_1162[19];
  assign _zz_1183 = _zz_1162[20];
  assign _zz_1184 = _zz_1162[21];
  assign _zz_1185 = _zz_1162[22];
  assign _zz_1186 = _zz_1162[23];
  assign _zz_1187 = _zz_1162[24];
  assign _zz_1188 = _zz_1162[25];
  assign _zz_1189 = _zz_1162[26];
  assign _zz_1190 = _zz_1162[27];
  assign _zz_1191 = _zz_1162[28];
  assign _zz_1192 = _zz_1162[29];
  assign _zz_1193 = _zz_1162[30];
  assign _zz_1194 = _zz_1162[31];
  assign _zz_1195 = _zz_1162[32];
  assign _zz_1196 = _zz_1162[33];
  assign _zz_1197 = _zz_1162[34];
  assign _zz_1198 = _zz_1162[35];
  assign _zz_1199 = _zz_1162[36];
  assign _zz_1200 = _zz_1162[37];
  assign _zz_1201 = _zz_1162[38];
  assign _zz_1202 = _zz_1162[39];
  assign _zz_1203 = _zz_1162[40];
  assign _zz_1204 = _zz_1162[41];
  assign _zz_1205 = _zz_1162[42];
  assign _zz_1206 = _zz_1162[43];
  assign _zz_1207 = _zz_1162[44];
  assign _zz_1208 = _zz_1162[45];
  assign _zz_1209 = _zz_1162[46];
  assign _zz_1210 = _zz_1162[47];
  assign _zz_1211 = _zz_1162[48];
  assign _zz_1212 = _zz_1162[49];
  assign _zz_1213 = _zz_1162[50];
  assign _zz_1214 = _zz_1162[51];
  assign _zz_1215 = _zz_1162[52];
  assign _zz_1216 = _zz_1162[53];
  assign _zz_1217 = _zz_1162[54];
  assign _zz_1218 = _zz_1162[55];
  assign _zz_1219 = _zz_1162[56];
  assign _zz_1220 = _zz_1162[57];
  assign _zz_1221 = _zz_1162[58];
  assign _zz_1222 = _zz_1162[59];
  assign _zz_1223 = _zz_1162[60];
  assign _zz_1224 = _zz_1162[61];
  assign _zz_1225 = _zz_1162[62];
  assign _zz_1226 = _zz_1162[63];
  assign _zz_1227 = _zz_1162[64];
  assign _zz_1228 = _zz_1162[65];
  assign _zz_1229 = _zz_1162[66];
  assign _zz_1230 = _zz_1162[67];
  assign _zz_1231 = _zz_1162[68];
  assign _zz_1232 = _zz_1162[69];
  assign _zz_1233 = _zz_1162[70];
  assign _zz_1234 = _zz_1162[71];
  assign _zz_1235 = _zz_1162[72];
  assign _zz_1236 = _zz_1162[73];
  assign _zz_1237 = _zz_1162[74];
  assign _zz_1238 = _zz_1162[75];
  assign _zz_1239 = _zz_1162[76];
  assign _zz_1240 = _zz_1162[77];
  assign _zz_1241 = _zz_1162[78];
  assign _zz_1242 = _zz_1162[79];
  assign _zz_1243 = _zz_1162[80];
  assign _zz_1244 = _zz_1162[81];
  assign _zz_1245 = _zz_1162[82];
  assign _zz_1246 = _zz_1162[83];
  assign _zz_1247 = _zz_1162[84];
  assign _zz_1248 = _zz_1162[85];
  assign _zz_1249 = _zz_1162[86];
  assign _zz_1250 = _zz_1162[87];
  assign _zz_1251 = _zz_1162[88];
  assign _zz_1252 = _zz_1162[89];
  assign _zz_1253 = _zz_1162[90];
  assign _zz_1254 = _zz_1162[91];
  assign _zz_1255 = _zz_1162[92];
  assign _zz_1256 = _zz_1162[93];
  assign _zz_1257 = _zz_1162[94];
  assign _zz_1258 = _zz_1162[95];
  assign _zz_1259 = _zz_1162[96];
  assign _zz_1260 = _zz_1162[97];
  assign _zz_1261 = _zz_1162[98];
  assign _zz_1262 = _zz_1162[99];
  assign _zz_1263 = _zz_1162[100];
  assign _zz_1264 = _zz_1162[101];
  assign _zz_1265 = _zz_1162[102];
  assign _zz_1266 = _zz_1162[103];
  assign _zz_1267 = _zz_1162[104];
  assign _zz_1268 = _zz_1162[105];
  assign _zz_1269 = _zz_1162[106];
  assign _zz_1270 = _zz_1162[107];
  assign _zz_1271 = _zz_1162[108];
  assign _zz_1272 = _zz_1162[109];
  assign _zz_1273 = _zz_1162[110];
  assign _zz_1274 = _zz_1162[111];
  assign _zz_1275 = _zz_1162[112];
  assign _zz_1276 = _zz_1162[113];
  assign _zz_1277 = _zz_1162[114];
  assign _zz_1278 = _zz_1162[115];
  assign _zz_1279 = _zz_1162[116];
  assign _zz_1280 = _zz_1162[117];
  assign _zz_1281 = _zz_1162[118];
  assign _zz_1282 = _zz_1162[119];
  assign _zz_1283 = _zz_1162[120];
  assign _zz_1284 = _zz_1162[121];
  assign _zz_1285 = _zz_1162[122];
  assign _zz_1286 = _zz_1162[123];
  assign _zz_1287 = _zz_1162[124];
  assign _zz_1288 = _zz_1162[125];
  assign _zz_1289 = _zz_1162[126];
  assign _zz_1290 = _zz_1162[127];
  assign cache_tag_3 = _zz_cache_tag_3;
  assign cache_hit_3 = ((cache_tag_3 == cpu_tag) && _zz_cache_hit_3);
  assign cache_mru_3 = _zz_cache_mru_3;
  assign _zz_1291 = ({127'd0,1'b1} <<< cpu_set_d1);
  assign _zz_1292 = _zz_1291[0];
  assign _zz_1293 = _zz_1291[1];
  assign _zz_1294 = _zz_1291[2];
  assign _zz_1295 = _zz_1291[3];
  assign _zz_1296 = _zz_1291[4];
  assign _zz_1297 = _zz_1291[5];
  assign _zz_1298 = _zz_1291[6];
  assign _zz_1299 = _zz_1291[7];
  assign _zz_1300 = _zz_1291[8];
  assign _zz_1301 = _zz_1291[9];
  assign _zz_1302 = _zz_1291[10];
  assign _zz_1303 = _zz_1291[11];
  assign _zz_1304 = _zz_1291[12];
  assign _zz_1305 = _zz_1291[13];
  assign _zz_1306 = _zz_1291[14];
  assign _zz_1307 = _zz_1291[15];
  assign _zz_1308 = _zz_1291[16];
  assign _zz_1309 = _zz_1291[17];
  assign _zz_1310 = _zz_1291[18];
  assign _zz_1311 = _zz_1291[19];
  assign _zz_1312 = _zz_1291[20];
  assign _zz_1313 = _zz_1291[21];
  assign _zz_1314 = _zz_1291[22];
  assign _zz_1315 = _zz_1291[23];
  assign _zz_1316 = _zz_1291[24];
  assign _zz_1317 = _zz_1291[25];
  assign _zz_1318 = _zz_1291[26];
  assign _zz_1319 = _zz_1291[27];
  assign _zz_1320 = _zz_1291[28];
  assign _zz_1321 = _zz_1291[29];
  assign _zz_1322 = _zz_1291[30];
  assign _zz_1323 = _zz_1291[31];
  assign _zz_1324 = _zz_1291[32];
  assign _zz_1325 = _zz_1291[33];
  assign _zz_1326 = _zz_1291[34];
  assign _zz_1327 = _zz_1291[35];
  assign _zz_1328 = _zz_1291[36];
  assign _zz_1329 = _zz_1291[37];
  assign _zz_1330 = _zz_1291[38];
  assign _zz_1331 = _zz_1291[39];
  assign _zz_1332 = _zz_1291[40];
  assign _zz_1333 = _zz_1291[41];
  assign _zz_1334 = _zz_1291[42];
  assign _zz_1335 = _zz_1291[43];
  assign _zz_1336 = _zz_1291[44];
  assign _zz_1337 = _zz_1291[45];
  assign _zz_1338 = _zz_1291[46];
  assign _zz_1339 = _zz_1291[47];
  assign _zz_1340 = _zz_1291[48];
  assign _zz_1341 = _zz_1291[49];
  assign _zz_1342 = _zz_1291[50];
  assign _zz_1343 = _zz_1291[51];
  assign _zz_1344 = _zz_1291[52];
  assign _zz_1345 = _zz_1291[53];
  assign _zz_1346 = _zz_1291[54];
  assign _zz_1347 = _zz_1291[55];
  assign _zz_1348 = _zz_1291[56];
  assign _zz_1349 = _zz_1291[57];
  assign _zz_1350 = _zz_1291[58];
  assign _zz_1351 = _zz_1291[59];
  assign _zz_1352 = _zz_1291[60];
  assign _zz_1353 = _zz_1291[61];
  assign _zz_1354 = _zz_1291[62];
  assign _zz_1355 = _zz_1291[63];
  assign _zz_1356 = _zz_1291[64];
  assign _zz_1357 = _zz_1291[65];
  assign _zz_1358 = _zz_1291[66];
  assign _zz_1359 = _zz_1291[67];
  assign _zz_1360 = _zz_1291[68];
  assign _zz_1361 = _zz_1291[69];
  assign _zz_1362 = _zz_1291[70];
  assign _zz_1363 = _zz_1291[71];
  assign _zz_1364 = _zz_1291[72];
  assign _zz_1365 = _zz_1291[73];
  assign _zz_1366 = _zz_1291[74];
  assign _zz_1367 = _zz_1291[75];
  assign _zz_1368 = _zz_1291[76];
  assign _zz_1369 = _zz_1291[77];
  assign _zz_1370 = _zz_1291[78];
  assign _zz_1371 = _zz_1291[79];
  assign _zz_1372 = _zz_1291[80];
  assign _zz_1373 = _zz_1291[81];
  assign _zz_1374 = _zz_1291[82];
  assign _zz_1375 = _zz_1291[83];
  assign _zz_1376 = _zz_1291[84];
  assign _zz_1377 = _zz_1291[85];
  assign _zz_1378 = _zz_1291[86];
  assign _zz_1379 = _zz_1291[87];
  assign _zz_1380 = _zz_1291[88];
  assign _zz_1381 = _zz_1291[89];
  assign _zz_1382 = _zz_1291[90];
  assign _zz_1383 = _zz_1291[91];
  assign _zz_1384 = _zz_1291[92];
  assign _zz_1385 = _zz_1291[93];
  assign _zz_1386 = _zz_1291[94];
  assign _zz_1387 = _zz_1291[95];
  assign _zz_1388 = _zz_1291[96];
  assign _zz_1389 = _zz_1291[97];
  assign _zz_1390 = _zz_1291[98];
  assign _zz_1391 = _zz_1291[99];
  assign _zz_1392 = _zz_1291[100];
  assign _zz_1393 = _zz_1291[101];
  assign _zz_1394 = _zz_1291[102];
  assign _zz_1395 = _zz_1291[103];
  assign _zz_1396 = _zz_1291[104];
  assign _zz_1397 = _zz_1291[105];
  assign _zz_1398 = _zz_1291[106];
  assign _zz_1399 = _zz_1291[107];
  assign _zz_1400 = _zz_1291[108];
  assign _zz_1401 = _zz_1291[109];
  assign _zz_1402 = _zz_1291[110];
  assign _zz_1403 = _zz_1291[111];
  assign _zz_1404 = _zz_1291[112];
  assign _zz_1405 = _zz_1291[113];
  assign _zz_1406 = _zz_1291[114];
  assign _zz_1407 = _zz_1291[115];
  assign _zz_1408 = _zz_1291[116];
  assign _zz_1409 = _zz_1291[117];
  assign _zz_1410 = _zz_1291[118];
  assign _zz_1411 = _zz_1291[119];
  assign _zz_1412 = _zz_1291[120];
  assign _zz_1413 = _zz_1291[121];
  assign _zz_1414 = _zz_1291[122];
  assign _zz_1415 = _zz_1291[123];
  assign _zz_1416 = _zz_1291[124];
  assign _zz_1417 = _zz_1291[125];
  assign _zz_1418 = _zz_1291[126];
  assign _zz_1419 = _zz_1291[127];
  assign cache_invld_d1_3 = (! _zz_cache_invld_d1_3);
  assign cache_lru_d1_3 = (! _zz_cache_lru_d1_3);
  assign cache_victim_3 = (cache_invld_d1_3 && cache_lru_d1_3);
  assign sram_banks_data_3 = sram_3_ports_rsp_payload_data;
  assign sram_banks_valid_3 = sram_3_ports_rsp_valid;
  assign when_ICache_l174_3 = (is_hit && (2'b11 == hit_id));
  always @(*) begin
    if(when_ICache_l174_3) begin
      sram_3_ports_cmd_payload_addr = cpu_bank_addr;
    end else begin
      if(when_ICache_l181_3) begin
        sram_3_ports_cmd_payload_addr = cpu_bank_addr_d1;
      end else begin
        if(when_ICache_l188_3) begin
          sram_3_ports_cmd_payload_addr = next_level_bank_addr;
        end else begin
          sram_3_ports_cmd_payload_addr = 7'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l174_3) begin
      sram_3_ports_cmd_valid = 1'b1;
    end else begin
      if(when_ICache_l181_3) begin
        sram_3_ports_cmd_valid = 1'b1;
      end else begin
        if(when_ICache_l188_3) begin
          sram_3_ports_cmd_valid = 1'b1;
        end else begin
          sram_3_ports_cmd_valid = 1'b0;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l174_3) begin
      sram_3_ports_cmd_payload_wen = 16'h0;
    end else begin
      if(when_ICache_l181_3) begin
        sram_3_ports_cmd_payload_wen = 16'h0;
      end else begin
        if(when_ICache_l188_3) begin
          sram_3_ports_cmd_payload_wen = (_zz_sram_3_ports_cmd_payload_wen <<< _zz_sram_3_ports_cmd_payload_wen_1);
        end else begin
          sram_3_ports_cmd_payload_wen = 16'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l174_3) begin
      sram_3_ports_cmd_payload_wdata = 512'h0;
    end else begin
      if(when_ICache_l181_3) begin
        sram_3_ports_cmd_payload_wdata = 512'h0;
      end else begin
        if(when_ICache_l188_3) begin
          sram_3_ports_cmd_payload_wdata = ({448'h0,next_level_rsp_payload_data} <<< _zz_sram_3_ports_cmd_payload_wdata);
        end else begin
          sram_3_ports_cmd_payload_wdata = 512'h0;
        end
      end
    end
  end

  always @(*) begin
    if(when_ICache_l174_3) begin
      sram_3_ports_cmd_payload_wstrb = 64'h0;
    end else begin
      if(when_ICache_l181_3) begin
        sram_3_ports_cmd_payload_wstrb = 64'h0;
      end else begin
        if(when_ICache_l188_3) begin
          sram_3_ports_cmd_payload_wstrb = ({56'h0,8'hff} <<< _zz_sram_3_ports_cmd_payload_wstrb);
        end else begin
          sram_3_ports_cmd_payload_wstrb = 64'h0;
        end
      end
    end
  end

  assign _zz_1552 = zz__zz_sram_3_ports_cmd_payload_wen(1'b0);
  always @(*) _zz_sram_3_ports_cmd_payload_wen = _zz_1552;
  assign when_ICache_l181_3 = (next_level_done && (2'b11 == evict_id_miss));
  assign when_ICache_l188_3 = (next_level_rsp_valid && (2'b11 == evict_id_miss));
  assign _zz_1420 = ({127'd0,1'b1} <<< flush_cnt_value);
  assign _zz_1421 = _zz_1420[0];
  assign _zz_1422 = _zz_1420[1];
  assign _zz_1423 = _zz_1420[2];
  assign _zz_1424 = _zz_1420[3];
  assign _zz_1425 = _zz_1420[4];
  assign _zz_1426 = _zz_1420[5];
  assign _zz_1427 = _zz_1420[6];
  assign _zz_1428 = _zz_1420[7];
  assign _zz_1429 = _zz_1420[8];
  assign _zz_1430 = _zz_1420[9];
  assign _zz_1431 = _zz_1420[10];
  assign _zz_1432 = _zz_1420[11];
  assign _zz_1433 = _zz_1420[12];
  assign _zz_1434 = _zz_1420[13];
  assign _zz_1435 = _zz_1420[14];
  assign _zz_1436 = _zz_1420[15];
  assign _zz_1437 = _zz_1420[16];
  assign _zz_1438 = _zz_1420[17];
  assign _zz_1439 = _zz_1420[18];
  assign _zz_1440 = _zz_1420[19];
  assign _zz_1441 = _zz_1420[20];
  assign _zz_1442 = _zz_1420[21];
  assign _zz_1443 = _zz_1420[22];
  assign _zz_1444 = _zz_1420[23];
  assign _zz_1445 = _zz_1420[24];
  assign _zz_1446 = _zz_1420[25];
  assign _zz_1447 = _zz_1420[26];
  assign _zz_1448 = _zz_1420[27];
  assign _zz_1449 = _zz_1420[28];
  assign _zz_1450 = _zz_1420[29];
  assign _zz_1451 = _zz_1420[30];
  assign _zz_1452 = _zz_1420[31];
  assign _zz_1453 = _zz_1420[32];
  assign _zz_1454 = _zz_1420[33];
  assign _zz_1455 = _zz_1420[34];
  assign _zz_1456 = _zz_1420[35];
  assign _zz_1457 = _zz_1420[36];
  assign _zz_1458 = _zz_1420[37];
  assign _zz_1459 = _zz_1420[38];
  assign _zz_1460 = _zz_1420[39];
  assign _zz_1461 = _zz_1420[40];
  assign _zz_1462 = _zz_1420[41];
  assign _zz_1463 = _zz_1420[42];
  assign _zz_1464 = _zz_1420[43];
  assign _zz_1465 = _zz_1420[44];
  assign _zz_1466 = _zz_1420[45];
  assign _zz_1467 = _zz_1420[46];
  assign _zz_1468 = _zz_1420[47];
  assign _zz_1469 = _zz_1420[48];
  assign _zz_1470 = _zz_1420[49];
  assign _zz_1471 = _zz_1420[50];
  assign _zz_1472 = _zz_1420[51];
  assign _zz_1473 = _zz_1420[52];
  assign _zz_1474 = _zz_1420[53];
  assign _zz_1475 = _zz_1420[54];
  assign _zz_1476 = _zz_1420[55];
  assign _zz_1477 = _zz_1420[56];
  assign _zz_1478 = _zz_1420[57];
  assign _zz_1479 = _zz_1420[58];
  assign _zz_1480 = _zz_1420[59];
  assign _zz_1481 = _zz_1420[60];
  assign _zz_1482 = _zz_1420[61];
  assign _zz_1483 = _zz_1420[62];
  assign _zz_1484 = _zz_1420[63];
  assign _zz_1485 = _zz_1420[64];
  assign _zz_1486 = _zz_1420[65];
  assign _zz_1487 = _zz_1420[66];
  assign _zz_1488 = _zz_1420[67];
  assign _zz_1489 = _zz_1420[68];
  assign _zz_1490 = _zz_1420[69];
  assign _zz_1491 = _zz_1420[70];
  assign _zz_1492 = _zz_1420[71];
  assign _zz_1493 = _zz_1420[72];
  assign _zz_1494 = _zz_1420[73];
  assign _zz_1495 = _zz_1420[74];
  assign _zz_1496 = _zz_1420[75];
  assign _zz_1497 = _zz_1420[76];
  assign _zz_1498 = _zz_1420[77];
  assign _zz_1499 = _zz_1420[78];
  assign _zz_1500 = _zz_1420[79];
  assign _zz_1501 = _zz_1420[80];
  assign _zz_1502 = _zz_1420[81];
  assign _zz_1503 = _zz_1420[82];
  assign _zz_1504 = _zz_1420[83];
  assign _zz_1505 = _zz_1420[84];
  assign _zz_1506 = _zz_1420[85];
  assign _zz_1507 = _zz_1420[86];
  assign _zz_1508 = _zz_1420[87];
  assign _zz_1509 = _zz_1420[88];
  assign _zz_1510 = _zz_1420[89];
  assign _zz_1511 = _zz_1420[90];
  assign _zz_1512 = _zz_1420[91];
  assign _zz_1513 = _zz_1420[92];
  assign _zz_1514 = _zz_1420[93];
  assign _zz_1515 = _zz_1420[94];
  assign _zz_1516 = _zz_1420[95];
  assign _zz_1517 = _zz_1420[96];
  assign _zz_1518 = _zz_1420[97];
  assign _zz_1519 = _zz_1420[98];
  assign _zz_1520 = _zz_1420[99];
  assign _zz_1521 = _zz_1420[100];
  assign _zz_1522 = _zz_1420[101];
  assign _zz_1523 = _zz_1420[102];
  assign _zz_1524 = _zz_1420[103];
  assign _zz_1525 = _zz_1420[104];
  assign _zz_1526 = _zz_1420[105];
  assign _zz_1527 = _zz_1420[106];
  assign _zz_1528 = _zz_1420[107];
  assign _zz_1529 = _zz_1420[108];
  assign _zz_1530 = _zz_1420[109];
  assign _zz_1531 = _zz_1420[110];
  assign _zz_1532 = _zz_1420[111];
  assign _zz_1533 = _zz_1420[112];
  assign _zz_1534 = _zz_1420[113];
  assign _zz_1535 = _zz_1420[114];
  assign _zz_1536 = _zz_1420[115];
  assign _zz_1537 = _zz_1420[116];
  assign _zz_1538 = _zz_1420[117];
  assign _zz_1539 = _zz_1420[118];
  assign _zz_1540 = _zz_1420[119];
  assign _zz_1541 = _zz_1420[120];
  assign _zz_1542 = _zz_1420[121];
  assign _zz_1543 = _zz_1420[122];
  assign _zz_1544 = _zz_1420[123];
  assign _zz_1545 = _zz_1420[124];
  assign _zz_1546 = _zz_1420[125];
  assign _zz_1547 = _zz_1420[126];
  assign _zz_1548 = _zz_1420[127];
  assign when_ICache_l210_3 = (is_hit && mru_full);
  assign when_ICache_l217_3 = (is_hit && cache_hit_3);
  assign when_ICache_l220_3 = (next_level_done && (2'b11 == evict_id_miss));
  assign when_ICache_l225_3 = (next_level_done && (2'b11 == evict_id_miss));
  assign when_ICache_l230_3 = (flush || is_miss);
  assign when_ICache_l233_3 = (flush_done || next_level_done);
  assign _zz_cpu_rsp_payload_data = _zz__zz_cpu_rsp_payload_data;
  assign _zz_cpu_rsp_payload_data_1 = _zz__zz_cpu_rsp_payload_data_1;
  assign cpu_rsp_payload_data = (is_hit_d1 ? _zz_cpu_rsp_payload_data_2 : _zz_cpu_rsp_payload_data_3);
  assign cpu_rsp_valid = (is_hit_d1 ? _zz_cpu_rsp_valid : _zz_cpu_rsp_valid_1);
  assign cpu_cmd_ready = cpu_cmd_ready_1;
  assign next_level_cmd_payload_addr = {cpu_addr_d1[63 : 6],6'h0};
  assign next_level_cmd_payload_len = 4'b0111;
  assign next_level_cmd_payload_size = 3'b011;
  assign next_level_cmd_valid = next_level_cmd_valid_1;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      ways_0_metas_0_vld <= 1'b0;
      ways_0_metas_0_tag <= 51'h0;
      ways_0_metas_0_mru <= 1'b0;
      ways_0_metas_1_vld <= 1'b0;
      ways_0_metas_1_tag <= 51'h0;
      ways_0_metas_1_mru <= 1'b0;
      ways_0_metas_2_vld <= 1'b0;
      ways_0_metas_2_tag <= 51'h0;
      ways_0_metas_2_mru <= 1'b0;
      ways_0_metas_3_vld <= 1'b0;
      ways_0_metas_3_tag <= 51'h0;
      ways_0_metas_3_mru <= 1'b0;
      ways_0_metas_4_vld <= 1'b0;
      ways_0_metas_4_tag <= 51'h0;
      ways_0_metas_4_mru <= 1'b0;
      ways_0_metas_5_vld <= 1'b0;
      ways_0_metas_5_tag <= 51'h0;
      ways_0_metas_5_mru <= 1'b0;
      ways_0_metas_6_vld <= 1'b0;
      ways_0_metas_6_tag <= 51'h0;
      ways_0_metas_6_mru <= 1'b0;
      ways_0_metas_7_vld <= 1'b0;
      ways_0_metas_7_tag <= 51'h0;
      ways_0_metas_7_mru <= 1'b0;
      ways_0_metas_8_vld <= 1'b0;
      ways_0_metas_8_tag <= 51'h0;
      ways_0_metas_8_mru <= 1'b0;
      ways_0_metas_9_vld <= 1'b0;
      ways_0_metas_9_tag <= 51'h0;
      ways_0_metas_9_mru <= 1'b0;
      ways_0_metas_10_vld <= 1'b0;
      ways_0_metas_10_tag <= 51'h0;
      ways_0_metas_10_mru <= 1'b0;
      ways_0_metas_11_vld <= 1'b0;
      ways_0_metas_11_tag <= 51'h0;
      ways_0_metas_11_mru <= 1'b0;
      ways_0_metas_12_vld <= 1'b0;
      ways_0_metas_12_tag <= 51'h0;
      ways_0_metas_12_mru <= 1'b0;
      ways_0_metas_13_vld <= 1'b0;
      ways_0_metas_13_tag <= 51'h0;
      ways_0_metas_13_mru <= 1'b0;
      ways_0_metas_14_vld <= 1'b0;
      ways_0_metas_14_tag <= 51'h0;
      ways_0_metas_14_mru <= 1'b0;
      ways_0_metas_15_vld <= 1'b0;
      ways_0_metas_15_tag <= 51'h0;
      ways_0_metas_15_mru <= 1'b0;
      ways_0_metas_16_vld <= 1'b0;
      ways_0_metas_16_tag <= 51'h0;
      ways_0_metas_16_mru <= 1'b0;
      ways_0_metas_17_vld <= 1'b0;
      ways_0_metas_17_tag <= 51'h0;
      ways_0_metas_17_mru <= 1'b0;
      ways_0_metas_18_vld <= 1'b0;
      ways_0_metas_18_tag <= 51'h0;
      ways_0_metas_18_mru <= 1'b0;
      ways_0_metas_19_vld <= 1'b0;
      ways_0_metas_19_tag <= 51'h0;
      ways_0_metas_19_mru <= 1'b0;
      ways_0_metas_20_vld <= 1'b0;
      ways_0_metas_20_tag <= 51'h0;
      ways_0_metas_20_mru <= 1'b0;
      ways_0_metas_21_vld <= 1'b0;
      ways_0_metas_21_tag <= 51'h0;
      ways_0_metas_21_mru <= 1'b0;
      ways_0_metas_22_vld <= 1'b0;
      ways_0_metas_22_tag <= 51'h0;
      ways_0_metas_22_mru <= 1'b0;
      ways_0_metas_23_vld <= 1'b0;
      ways_0_metas_23_tag <= 51'h0;
      ways_0_metas_23_mru <= 1'b0;
      ways_0_metas_24_vld <= 1'b0;
      ways_0_metas_24_tag <= 51'h0;
      ways_0_metas_24_mru <= 1'b0;
      ways_0_metas_25_vld <= 1'b0;
      ways_0_metas_25_tag <= 51'h0;
      ways_0_metas_25_mru <= 1'b0;
      ways_0_metas_26_vld <= 1'b0;
      ways_0_metas_26_tag <= 51'h0;
      ways_0_metas_26_mru <= 1'b0;
      ways_0_metas_27_vld <= 1'b0;
      ways_0_metas_27_tag <= 51'h0;
      ways_0_metas_27_mru <= 1'b0;
      ways_0_metas_28_vld <= 1'b0;
      ways_0_metas_28_tag <= 51'h0;
      ways_0_metas_28_mru <= 1'b0;
      ways_0_metas_29_vld <= 1'b0;
      ways_0_metas_29_tag <= 51'h0;
      ways_0_metas_29_mru <= 1'b0;
      ways_0_metas_30_vld <= 1'b0;
      ways_0_metas_30_tag <= 51'h0;
      ways_0_metas_30_mru <= 1'b0;
      ways_0_metas_31_vld <= 1'b0;
      ways_0_metas_31_tag <= 51'h0;
      ways_0_metas_31_mru <= 1'b0;
      ways_0_metas_32_vld <= 1'b0;
      ways_0_metas_32_tag <= 51'h0;
      ways_0_metas_32_mru <= 1'b0;
      ways_0_metas_33_vld <= 1'b0;
      ways_0_metas_33_tag <= 51'h0;
      ways_0_metas_33_mru <= 1'b0;
      ways_0_metas_34_vld <= 1'b0;
      ways_0_metas_34_tag <= 51'h0;
      ways_0_metas_34_mru <= 1'b0;
      ways_0_metas_35_vld <= 1'b0;
      ways_0_metas_35_tag <= 51'h0;
      ways_0_metas_35_mru <= 1'b0;
      ways_0_metas_36_vld <= 1'b0;
      ways_0_metas_36_tag <= 51'h0;
      ways_0_metas_36_mru <= 1'b0;
      ways_0_metas_37_vld <= 1'b0;
      ways_0_metas_37_tag <= 51'h0;
      ways_0_metas_37_mru <= 1'b0;
      ways_0_metas_38_vld <= 1'b0;
      ways_0_metas_38_tag <= 51'h0;
      ways_0_metas_38_mru <= 1'b0;
      ways_0_metas_39_vld <= 1'b0;
      ways_0_metas_39_tag <= 51'h0;
      ways_0_metas_39_mru <= 1'b0;
      ways_0_metas_40_vld <= 1'b0;
      ways_0_metas_40_tag <= 51'h0;
      ways_0_metas_40_mru <= 1'b0;
      ways_0_metas_41_vld <= 1'b0;
      ways_0_metas_41_tag <= 51'h0;
      ways_0_metas_41_mru <= 1'b0;
      ways_0_metas_42_vld <= 1'b0;
      ways_0_metas_42_tag <= 51'h0;
      ways_0_metas_42_mru <= 1'b0;
      ways_0_metas_43_vld <= 1'b0;
      ways_0_metas_43_tag <= 51'h0;
      ways_0_metas_43_mru <= 1'b0;
      ways_0_metas_44_vld <= 1'b0;
      ways_0_metas_44_tag <= 51'h0;
      ways_0_metas_44_mru <= 1'b0;
      ways_0_metas_45_vld <= 1'b0;
      ways_0_metas_45_tag <= 51'h0;
      ways_0_metas_45_mru <= 1'b0;
      ways_0_metas_46_vld <= 1'b0;
      ways_0_metas_46_tag <= 51'h0;
      ways_0_metas_46_mru <= 1'b0;
      ways_0_metas_47_vld <= 1'b0;
      ways_0_metas_47_tag <= 51'h0;
      ways_0_metas_47_mru <= 1'b0;
      ways_0_metas_48_vld <= 1'b0;
      ways_0_metas_48_tag <= 51'h0;
      ways_0_metas_48_mru <= 1'b0;
      ways_0_metas_49_vld <= 1'b0;
      ways_0_metas_49_tag <= 51'h0;
      ways_0_metas_49_mru <= 1'b0;
      ways_0_metas_50_vld <= 1'b0;
      ways_0_metas_50_tag <= 51'h0;
      ways_0_metas_50_mru <= 1'b0;
      ways_0_metas_51_vld <= 1'b0;
      ways_0_metas_51_tag <= 51'h0;
      ways_0_metas_51_mru <= 1'b0;
      ways_0_metas_52_vld <= 1'b0;
      ways_0_metas_52_tag <= 51'h0;
      ways_0_metas_52_mru <= 1'b0;
      ways_0_metas_53_vld <= 1'b0;
      ways_0_metas_53_tag <= 51'h0;
      ways_0_metas_53_mru <= 1'b0;
      ways_0_metas_54_vld <= 1'b0;
      ways_0_metas_54_tag <= 51'h0;
      ways_0_metas_54_mru <= 1'b0;
      ways_0_metas_55_vld <= 1'b0;
      ways_0_metas_55_tag <= 51'h0;
      ways_0_metas_55_mru <= 1'b0;
      ways_0_metas_56_vld <= 1'b0;
      ways_0_metas_56_tag <= 51'h0;
      ways_0_metas_56_mru <= 1'b0;
      ways_0_metas_57_vld <= 1'b0;
      ways_0_metas_57_tag <= 51'h0;
      ways_0_metas_57_mru <= 1'b0;
      ways_0_metas_58_vld <= 1'b0;
      ways_0_metas_58_tag <= 51'h0;
      ways_0_metas_58_mru <= 1'b0;
      ways_0_metas_59_vld <= 1'b0;
      ways_0_metas_59_tag <= 51'h0;
      ways_0_metas_59_mru <= 1'b0;
      ways_0_metas_60_vld <= 1'b0;
      ways_0_metas_60_tag <= 51'h0;
      ways_0_metas_60_mru <= 1'b0;
      ways_0_metas_61_vld <= 1'b0;
      ways_0_metas_61_tag <= 51'h0;
      ways_0_metas_61_mru <= 1'b0;
      ways_0_metas_62_vld <= 1'b0;
      ways_0_metas_62_tag <= 51'h0;
      ways_0_metas_62_mru <= 1'b0;
      ways_0_metas_63_vld <= 1'b0;
      ways_0_metas_63_tag <= 51'h0;
      ways_0_metas_63_mru <= 1'b0;
      ways_0_metas_64_vld <= 1'b0;
      ways_0_metas_64_tag <= 51'h0;
      ways_0_metas_64_mru <= 1'b0;
      ways_0_metas_65_vld <= 1'b0;
      ways_0_metas_65_tag <= 51'h0;
      ways_0_metas_65_mru <= 1'b0;
      ways_0_metas_66_vld <= 1'b0;
      ways_0_metas_66_tag <= 51'h0;
      ways_0_metas_66_mru <= 1'b0;
      ways_0_metas_67_vld <= 1'b0;
      ways_0_metas_67_tag <= 51'h0;
      ways_0_metas_67_mru <= 1'b0;
      ways_0_metas_68_vld <= 1'b0;
      ways_0_metas_68_tag <= 51'h0;
      ways_0_metas_68_mru <= 1'b0;
      ways_0_metas_69_vld <= 1'b0;
      ways_0_metas_69_tag <= 51'h0;
      ways_0_metas_69_mru <= 1'b0;
      ways_0_metas_70_vld <= 1'b0;
      ways_0_metas_70_tag <= 51'h0;
      ways_0_metas_70_mru <= 1'b0;
      ways_0_metas_71_vld <= 1'b0;
      ways_0_metas_71_tag <= 51'h0;
      ways_0_metas_71_mru <= 1'b0;
      ways_0_metas_72_vld <= 1'b0;
      ways_0_metas_72_tag <= 51'h0;
      ways_0_metas_72_mru <= 1'b0;
      ways_0_metas_73_vld <= 1'b0;
      ways_0_metas_73_tag <= 51'h0;
      ways_0_metas_73_mru <= 1'b0;
      ways_0_metas_74_vld <= 1'b0;
      ways_0_metas_74_tag <= 51'h0;
      ways_0_metas_74_mru <= 1'b0;
      ways_0_metas_75_vld <= 1'b0;
      ways_0_metas_75_tag <= 51'h0;
      ways_0_metas_75_mru <= 1'b0;
      ways_0_metas_76_vld <= 1'b0;
      ways_0_metas_76_tag <= 51'h0;
      ways_0_metas_76_mru <= 1'b0;
      ways_0_metas_77_vld <= 1'b0;
      ways_0_metas_77_tag <= 51'h0;
      ways_0_metas_77_mru <= 1'b0;
      ways_0_metas_78_vld <= 1'b0;
      ways_0_metas_78_tag <= 51'h0;
      ways_0_metas_78_mru <= 1'b0;
      ways_0_metas_79_vld <= 1'b0;
      ways_0_metas_79_tag <= 51'h0;
      ways_0_metas_79_mru <= 1'b0;
      ways_0_metas_80_vld <= 1'b0;
      ways_0_metas_80_tag <= 51'h0;
      ways_0_metas_80_mru <= 1'b0;
      ways_0_metas_81_vld <= 1'b0;
      ways_0_metas_81_tag <= 51'h0;
      ways_0_metas_81_mru <= 1'b0;
      ways_0_metas_82_vld <= 1'b0;
      ways_0_metas_82_tag <= 51'h0;
      ways_0_metas_82_mru <= 1'b0;
      ways_0_metas_83_vld <= 1'b0;
      ways_0_metas_83_tag <= 51'h0;
      ways_0_metas_83_mru <= 1'b0;
      ways_0_metas_84_vld <= 1'b0;
      ways_0_metas_84_tag <= 51'h0;
      ways_0_metas_84_mru <= 1'b0;
      ways_0_metas_85_vld <= 1'b0;
      ways_0_metas_85_tag <= 51'h0;
      ways_0_metas_85_mru <= 1'b0;
      ways_0_metas_86_vld <= 1'b0;
      ways_0_metas_86_tag <= 51'h0;
      ways_0_metas_86_mru <= 1'b0;
      ways_0_metas_87_vld <= 1'b0;
      ways_0_metas_87_tag <= 51'h0;
      ways_0_metas_87_mru <= 1'b0;
      ways_0_metas_88_vld <= 1'b0;
      ways_0_metas_88_tag <= 51'h0;
      ways_0_metas_88_mru <= 1'b0;
      ways_0_metas_89_vld <= 1'b0;
      ways_0_metas_89_tag <= 51'h0;
      ways_0_metas_89_mru <= 1'b0;
      ways_0_metas_90_vld <= 1'b0;
      ways_0_metas_90_tag <= 51'h0;
      ways_0_metas_90_mru <= 1'b0;
      ways_0_metas_91_vld <= 1'b0;
      ways_0_metas_91_tag <= 51'h0;
      ways_0_metas_91_mru <= 1'b0;
      ways_0_metas_92_vld <= 1'b0;
      ways_0_metas_92_tag <= 51'h0;
      ways_0_metas_92_mru <= 1'b0;
      ways_0_metas_93_vld <= 1'b0;
      ways_0_metas_93_tag <= 51'h0;
      ways_0_metas_93_mru <= 1'b0;
      ways_0_metas_94_vld <= 1'b0;
      ways_0_metas_94_tag <= 51'h0;
      ways_0_metas_94_mru <= 1'b0;
      ways_0_metas_95_vld <= 1'b0;
      ways_0_metas_95_tag <= 51'h0;
      ways_0_metas_95_mru <= 1'b0;
      ways_0_metas_96_vld <= 1'b0;
      ways_0_metas_96_tag <= 51'h0;
      ways_0_metas_96_mru <= 1'b0;
      ways_0_metas_97_vld <= 1'b0;
      ways_0_metas_97_tag <= 51'h0;
      ways_0_metas_97_mru <= 1'b0;
      ways_0_metas_98_vld <= 1'b0;
      ways_0_metas_98_tag <= 51'h0;
      ways_0_metas_98_mru <= 1'b0;
      ways_0_metas_99_vld <= 1'b0;
      ways_0_metas_99_tag <= 51'h0;
      ways_0_metas_99_mru <= 1'b0;
      ways_0_metas_100_vld <= 1'b0;
      ways_0_metas_100_tag <= 51'h0;
      ways_0_metas_100_mru <= 1'b0;
      ways_0_metas_101_vld <= 1'b0;
      ways_0_metas_101_tag <= 51'h0;
      ways_0_metas_101_mru <= 1'b0;
      ways_0_metas_102_vld <= 1'b0;
      ways_0_metas_102_tag <= 51'h0;
      ways_0_metas_102_mru <= 1'b0;
      ways_0_metas_103_vld <= 1'b0;
      ways_0_metas_103_tag <= 51'h0;
      ways_0_metas_103_mru <= 1'b0;
      ways_0_metas_104_vld <= 1'b0;
      ways_0_metas_104_tag <= 51'h0;
      ways_0_metas_104_mru <= 1'b0;
      ways_0_metas_105_vld <= 1'b0;
      ways_0_metas_105_tag <= 51'h0;
      ways_0_metas_105_mru <= 1'b0;
      ways_0_metas_106_vld <= 1'b0;
      ways_0_metas_106_tag <= 51'h0;
      ways_0_metas_106_mru <= 1'b0;
      ways_0_metas_107_vld <= 1'b0;
      ways_0_metas_107_tag <= 51'h0;
      ways_0_metas_107_mru <= 1'b0;
      ways_0_metas_108_vld <= 1'b0;
      ways_0_metas_108_tag <= 51'h0;
      ways_0_metas_108_mru <= 1'b0;
      ways_0_metas_109_vld <= 1'b0;
      ways_0_metas_109_tag <= 51'h0;
      ways_0_metas_109_mru <= 1'b0;
      ways_0_metas_110_vld <= 1'b0;
      ways_0_metas_110_tag <= 51'h0;
      ways_0_metas_110_mru <= 1'b0;
      ways_0_metas_111_vld <= 1'b0;
      ways_0_metas_111_tag <= 51'h0;
      ways_0_metas_111_mru <= 1'b0;
      ways_0_metas_112_vld <= 1'b0;
      ways_0_metas_112_tag <= 51'h0;
      ways_0_metas_112_mru <= 1'b0;
      ways_0_metas_113_vld <= 1'b0;
      ways_0_metas_113_tag <= 51'h0;
      ways_0_metas_113_mru <= 1'b0;
      ways_0_metas_114_vld <= 1'b0;
      ways_0_metas_114_tag <= 51'h0;
      ways_0_metas_114_mru <= 1'b0;
      ways_0_metas_115_vld <= 1'b0;
      ways_0_metas_115_tag <= 51'h0;
      ways_0_metas_115_mru <= 1'b0;
      ways_0_metas_116_vld <= 1'b0;
      ways_0_metas_116_tag <= 51'h0;
      ways_0_metas_116_mru <= 1'b0;
      ways_0_metas_117_vld <= 1'b0;
      ways_0_metas_117_tag <= 51'h0;
      ways_0_metas_117_mru <= 1'b0;
      ways_0_metas_118_vld <= 1'b0;
      ways_0_metas_118_tag <= 51'h0;
      ways_0_metas_118_mru <= 1'b0;
      ways_0_metas_119_vld <= 1'b0;
      ways_0_metas_119_tag <= 51'h0;
      ways_0_metas_119_mru <= 1'b0;
      ways_0_metas_120_vld <= 1'b0;
      ways_0_metas_120_tag <= 51'h0;
      ways_0_metas_120_mru <= 1'b0;
      ways_0_metas_121_vld <= 1'b0;
      ways_0_metas_121_tag <= 51'h0;
      ways_0_metas_121_mru <= 1'b0;
      ways_0_metas_122_vld <= 1'b0;
      ways_0_metas_122_tag <= 51'h0;
      ways_0_metas_122_mru <= 1'b0;
      ways_0_metas_123_vld <= 1'b0;
      ways_0_metas_123_tag <= 51'h0;
      ways_0_metas_123_mru <= 1'b0;
      ways_0_metas_124_vld <= 1'b0;
      ways_0_metas_124_tag <= 51'h0;
      ways_0_metas_124_mru <= 1'b0;
      ways_0_metas_125_vld <= 1'b0;
      ways_0_metas_125_tag <= 51'h0;
      ways_0_metas_125_mru <= 1'b0;
      ways_0_metas_126_vld <= 1'b0;
      ways_0_metas_126_tag <= 51'h0;
      ways_0_metas_126_mru <= 1'b0;
      ways_0_metas_127_vld <= 1'b0;
      ways_0_metas_127_tag <= 51'h0;
      ways_0_metas_127_mru <= 1'b0;
      ways_1_metas_0_vld <= 1'b0;
      ways_1_metas_0_tag <= 51'h0;
      ways_1_metas_0_mru <= 1'b0;
      ways_1_metas_1_vld <= 1'b0;
      ways_1_metas_1_tag <= 51'h0;
      ways_1_metas_1_mru <= 1'b0;
      ways_1_metas_2_vld <= 1'b0;
      ways_1_metas_2_tag <= 51'h0;
      ways_1_metas_2_mru <= 1'b0;
      ways_1_metas_3_vld <= 1'b0;
      ways_1_metas_3_tag <= 51'h0;
      ways_1_metas_3_mru <= 1'b0;
      ways_1_metas_4_vld <= 1'b0;
      ways_1_metas_4_tag <= 51'h0;
      ways_1_metas_4_mru <= 1'b0;
      ways_1_metas_5_vld <= 1'b0;
      ways_1_metas_5_tag <= 51'h0;
      ways_1_metas_5_mru <= 1'b0;
      ways_1_metas_6_vld <= 1'b0;
      ways_1_metas_6_tag <= 51'h0;
      ways_1_metas_6_mru <= 1'b0;
      ways_1_metas_7_vld <= 1'b0;
      ways_1_metas_7_tag <= 51'h0;
      ways_1_metas_7_mru <= 1'b0;
      ways_1_metas_8_vld <= 1'b0;
      ways_1_metas_8_tag <= 51'h0;
      ways_1_metas_8_mru <= 1'b0;
      ways_1_metas_9_vld <= 1'b0;
      ways_1_metas_9_tag <= 51'h0;
      ways_1_metas_9_mru <= 1'b0;
      ways_1_metas_10_vld <= 1'b0;
      ways_1_metas_10_tag <= 51'h0;
      ways_1_metas_10_mru <= 1'b0;
      ways_1_metas_11_vld <= 1'b0;
      ways_1_metas_11_tag <= 51'h0;
      ways_1_metas_11_mru <= 1'b0;
      ways_1_metas_12_vld <= 1'b0;
      ways_1_metas_12_tag <= 51'h0;
      ways_1_metas_12_mru <= 1'b0;
      ways_1_metas_13_vld <= 1'b0;
      ways_1_metas_13_tag <= 51'h0;
      ways_1_metas_13_mru <= 1'b0;
      ways_1_metas_14_vld <= 1'b0;
      ways_1_metas_14_tag <= 51'h0;
      ways_1_metas_14_mru <= 1'b0;
      ways_1_metas_15_vld <= 1'b0;
      ways_1_metas_15_tag <= 51'h0;
      ways_1_metas_15_mru <= 1'b0;
      ways_1_metas_16_vld <= 1'b0;
      ways_1_metas_16_tag <= 51'h0;
      ways_1_metas_16_mru <= 1'b0;
      ways_1_metas_17_vld <= 1'b0;
      ways_1_metas_17_tag <= 51'h0;
      ways_1_metas_17_mru <= 1'b0;
      ways_1_metas_18_vld <= 1'b0;
      ways_1_metas_18_tag <= 51'h0;
      ways_1_metas_18_mru <= 1'b0;
      ways_1_metas_19_vld <= 1'b0;
      ways_1_metas_19_tag <= 51'h0;
      ways_1_metas_19_mru <= 1'b0;
      ways_1_metas_20_vld <= 1'b0;
      ways_1_metas_20_tag <= 51'h0;
      ways_1_metas_20_mru <= 1'b0;
      ways_1_metas_21_vld <= 1'b0;
      ways_1_metas_21_tag <= 51'h0;
      ways_1_metas_21_mru <= 1'b0;
      ways_1_metas_22_vld <= 1'b0;
      ways_1_metas_22_tag <= 51'h0;
      ways_1_metas_22_mru <= 1'b0;
      ways_1_metas_23_vld <= 1'b0;
      ways_1_metas_23_tag <= 51'h0;
      ways_1_metas_23_mru <= 1'b0;
      ways_1_metas_24_vld <= 1'b0;
      ways_1_metas_24_tag <= 51'h0;
      ways_1_metas_24_mru <= 1'b0;
      ways_1_metas_25_vld <= 1'b0;
      ways_1_metas_25_tag <= 51'h0;
      ways_1_metas_25_mru <= 1'b0;
      ways_1_metas_26_vld <= 1'b0;
      ways_1_metas_26_tag <= 51'h0;
      ways_1_metas_26_mru <= 1'b0;
      ways_1_metas_27_vld <= 1'b0;
      ways_1_metas_27_tag <= 51'h0;
      ways_1_metas_27_mru <= 1'b0;
      ways_1_metas_28_vld <= 1'b0;
      ways_1_metas_28_tag <= 51'h0;
      ways_1_metas_28_mru <= 1'b0;
      ways_1_metas_29_vld <= 1'b0;
      ways_1_metas_29_tag <= 51'h0;
      ways_1_metas_29_mru <= 1'b0;
      ways_1_metas_30_vld <= 1'b0;
      ways_1_metas_30_tag <= 51'h0;
      ways_1_metas_30_mru <= 1'b0;
      ways_1_metas_31_vld <= 1'b0;
      ways_1_metas_31_tag <= 51'h0;
      ways_1_metas_31_mru <= 1'b0;
      ways_1_metas_32_vld <= 1'b0;
      ways_1_metas_32_tag <= 51'h0;
      ways_1_metas_32_mru <= 1'b0;
      ways_1_metas_33_vld <= 1'b0;
      ways_1_metas_33_tag <= 51'h0;
      ways_1_metas_33_mru <= 1'b0;
      ways_1_metas_34_vld <= 1'b0;
      ways_1_metas_34_tag <= 51'h0;
      ways_1_metas_34_mru <= 1'b0;
      ways_1_metas_35_vld <= 1'b0;
      ways_1_metas_35_tag <= 51'h0;
      ways_1_metas_35_mru <= 1'b0;
      ways_1_metas_36_vld <= 1'b0;
      ways_1_metas_36_tag <= 51'h0;
      ways_1_metas_36_mru <= 1'b0;
      ways_1_metas_37_vld <= 1'b0;
      ways_1_metas_37_tag <= 51'h0;
      ways_1_metas_37_mru <= 1'b0;
      ways_1_metas_38_vld <= 1'b0;
      ways_1_metas_38_tag <= 51'h0;
      ways_1_metas_38_mru <= 1'b0;
      ways_1_metas_39_vld <= 1'b0;
      ways_1_metas_39_tag <= 51'h0;
      ways_1_metas_39_mru <= 1'b0;
      ways_1_metas_40_vld <= 1'b0;
      ways_1_metas_40_tag <= 51'h0;
      ways_1_metas_40_mru <= 1'b0;
      ways_1_metas_41_vld <= 1'b0;
      ways_1_metas_41_tag <= 51'h0;
      ways_1_metas_41_mru <= 1'b0;
      ways_1_metas_42_vld <= 1'b0;
      ways_1_metas_42_tag <= 51'h0;
      ways_1_metas_42_mru <= 1'b0;
      ways_1_metas_43_vld <= 1'b0;
      ways_1_metas_43_tag <= 51'h0;
      ways_1_metas_43_mru <= 1'b0;
      ways_1_metas_44_vld <= 1'b0;
      ways_1_metas_44_tag <= 51'h0;
      ways_1_metas_44_mru <= 1'b0;
      ways_1_metas_45_vld <= 1'b0;
      ways_1_metas_45_tag <= 51'h0;
      ways_1_metas_45_mru <= 1'b0;
      ways_1_metas_46_vld <= 1'b0;
      ways_1_metas_46_tag <= 51'h0;
      ways_1_metas_46_mru <= 1'b0;
      ways_1_metas_47_vld <= 1'b0;
      ways_1_metas_47_tag <= 51'h0;
      ways_1_metas_47_mru <= 1'b0;
      ways_1_metas_48_vld <= 1'b0;
      ways_1_metas_48_tag <= 51'h0;
      ways_1_metas_48_mru <= 1'b0;
      ways_1_metas_49_vld <= 1'b0;
      ways_1_metas_49_tag <= 51'h0;
      ways_1_metas_49_mru <= 1'b0;
      ways_1_metas_50_vld <= 1'b0;
      ways_1_metas_50_tag <= 51'h0;
      ways_1_metas_50_mru <= 1'b0;
      ways_1_metas_51_vld <= 1'b0;
      ways_1_metas_51_tag <= 51'h0;
      ways_1_metas_51_mru <= 1'b0;
      ways_1_metas_52_vld <= 1'b0;
      ways_1_metas_52_tag <= 51'h0;
      ways_1_metas_52_mru <= 1'b0;
      ways_1_metas_53_vld <= 1'b0;
      ways_1_metas_53_tag <= 51'h0;
      ways_1_metas_53_mru <= 1'b0;
      ways_1_metas_54_vld <= 1'b0;
      ways_1_metas_54_tag <= 51'h0;
      ways_1_metas_54_mru <= 1'b0;
      ways_1_metas_55_vld <= 1'b0;
      ways_1_metas_55_tag <= 51'h0;
      ways_1_metas_55_mru <= 1'b0;
      ways_1_metas_56_vld <= 1'b0;
      ways_1_metas_56_tag <= 51'h0;
      ways_1_metas_56_mru <= 1'b0;
      ways_1_metas_57_vld <= 1'b0;
      ways_1_metas_57_tag <= 51'h0;
      ways_1_metas_57_mru <= 1'b0;
      ways_1_metas_58_vld <= 1'b0;
      ways_1_metas_58_tag <= 51'h0;
      ways_1_metas_58_mru <= 1'b0;
      ways_1_metas_59_vld <= 1'b0;
      ways_1_metas_59_tag <= 51'h0;
      ways_1_metas_59_mru <= 1'b0;
      ways_1_metas_60_vld <= 1'b0;
      ways_1_metas_60_tag <= 51'h0;
      ways_1_metas_60_mru <= 1'b0;
      ways_1_metas_61_vld <= 1'b0;
      ways_1_metas_61_tag <= 51'h0;
      ways_1_metas_61_mru <= 1'b0;
      ways_1_metas_62_vld <= 1'b0;
      ways_1_metas_62_tag <= 51'h0;
      ways_1_metas_62_mru <= 1'b0;
      ways_1_metas_63_vld <= 1'b0;
      ways_1_metas_63_tag <= 51'h0;
      ways_1_metas_63_mru <= 1'b0;
      ways_1_metas_64_vld <= 1'b0;
      ways_1_metas_64_tag <= 51'h0;
      ways_1_metas_64_mru <= 1'b0;
      ways_1_metas_65_vld <= 1'b0;
      ways_1_metas_65_tag <= 51'h0;
      ways_1_metas_65_mru <= 1'b0;
      ways_1_metas_66_vld <= 1'b0;
      ways_1_metas_66_tag <= 51'h0;
      ways_1_metas_66_mru <= 1'b0;
      ways_1_metas_67_vld <= 1'b0;
      ways_1_metas_67_tag <= 51'h0;
      ways_1_metas_67_mru <= 1'b0;
      ways_1_metas_68_vld <= 1'b0;
      ways_1_metas_68_tag <= 51'h0;
      ways_1_metas_68_mru <= 1'b0;
      ways_1_metas_69_vld <= 1'b0;
      ways_1_metas_69_tag <= 51'h0;
      ways_1_metas_69_mru <= 1'b0;
      ways_1_metas_70_vld <= 1'b0;
      ways_1_metas_70_tag <= 51'h0;
      ways_1_metas_70_mru <= 1'b0;
      ways_1_metas_71_vld <= 1'b0;
      ways_1_metas_71_tag <= 51'h0;
      ways_1_metas_71_mru <= 1'b0;
      ways_1_metas_72_vld <= 1'b0;
      ways_1_metas_72_tag <= 51'h0;
      ways_1_metas_72_mru <= 1'b0;
      ways_1_metas_73_vld <= 1'b0;
      ways_1_metas_73_tag <= 51'h0;
      ways_1_metas_73_mru <= 1'b0;
      ways_1_metas_74_vld <= 1'b0;
      ways_1_metas_74_tag <= 51'h0;
      ways_1_metas_74_mru <= 1'b0;
      ways_1_metas_75_vld <= 1'b0;
      ways_1_metas_75_tag <= 51'h0;
      ways_1_metas_75_mru <= 1'b0;
      ways_1_metas_76_vld <= 1'b0;
      ways_1_metas_76_tag <= 51'h0;
      ways_1_metas_76_mru <= 1'b0;
      ways_1_metas_77_vld <= 1'b0;
      ways_1_metas_77_tag <= 51'h0;
      ways_1_metas_77_mru <= 1'b0;
      ways_1_metas_78_vld <= 1'b0;
      ways_1_metas_78_tag <= 51'h0;
      ways_1_metas_78_mru <= 1'b0;
      ways_1_metas_79_vld <= 1'b0;
      ways_1_metas_79_tag <= 51'h0;
      ways_1_metas_79_mru <= 1'b0;
      ways_1_metas_80_vld <= 1'b0;
      ways_1_metas_80_tag <= 51'h0;
      ways_1_metas_80_mru <= 1'b0;
      ways_1_metas_81_vld <= 1'b0;
      ways_1_metas_81_tag <= 51'h0;
      ways_1_metas_81_mru <= 1'b0;
      ways_1_metas_82_vld <= 1'b0;
      ways_1_metas_82_tag <= 51'h0;
      ways_1_metas_82_mru <= 1'b0;
      ways_1_metas_83_vld <= 1'b0;
      ways_1_metas_83_tag <= 51'h0;
      ways_1_metas_83_mru <= 1'b0;
      ways_1_metas_84_vld <= 1'b0;
      ways_1_metas_84_tag <= 51'h0;
      ways_1_metas_84_mru <= 1'b0;
      ways_1_metas_85_vld <= 1'b0;
      ways_1_metas_85_tag <= 51'h0;
      ways_1_metas_85_mru <= 1'b0;
      ways_1_metas_86_vld <= 1'b0;
      ways_1_metas_86_tag <= 51'h0;
      ways_1_metas_86_mru <= 1'b0;
      ways_1_metas_87_vld <= 1'b0;
      ways_1_metas_87_tag <= 51'h0;
      ways_1_metas_87_mru <= 1'b0;
      ways_1_metas_88_vld <= 1'b0;
      ways_1_metas_88_tag <= 51'h0;
      ways_1_metas_88_mru <= 1'b0;
      ways_1_metas_89_vld <= 1'b0;
      ways_1_metas_89_tag <= 51'h0;
      ways_1_metas_89_mru <= 1'b0;
      ways_1_metas_90_vld <= 1'b0;
      ways_1_metas_90_tag <= 51'h0;
      ways_1_metas_90_mru <= 1'b0;
      ways_1_metas_91_vld <= 1'b0;
      ways_1_metas_91_tag <= 51'h0;
      ways_1_metas_91_mru <= 1'b0;
      ways_1_metas_92_vld <= 1'b0;
      ways_1_metas_92_tag <= 51'h0;
      ways_1_metas_92_mru <= 1'b0;
      ways_1_metas_93_vld <= 1'b0;
      ways_1_metas_93_tag <= 51'h0;
      ways_1_metas_93_mru <= 1'b0;
      ways_1_metas_94_vld <= 1'b0;
      ways_1_metas_94_tag <= 51'h0;
      ways_1_metas_94_mru <= 1'b0;
      ways_1_metas_95_vld <= 1'b0;
      ways_1_metas_95_tag <= 51'h0;
      ways_1_metas_95_mru <= 1'b0;
      ways_1_metas_96_vld <= 1'b0;
      ways_1_metas_96_tag <= 51'h0;
      ways_1_metas_96_mru <= 1'b0;
      ways_1_metas_97_vld <= 1'b0;
      ways_1_metas_97_tag <= 51'h0;
      ways_1_metas_97_mru <= 1'b0;
      ways_1_metas_98_vld <= 1'b0;
      ways_1_metas_98_tag <= 51'h0;
      ways_1_metas_98_mru <= 1'b0;
      ways_1_metas_99_vld <= 1'b0;
      ways_1_metas_99_tag <= 51'h0;
      ways_1_metas_99_mru <= 1'b0;
      ways_1_metas_100_vld <= 1'b0;
      ways_1_metas_100_tag <= 51'h0;
      ways_1_metas_100_mru <= 1'b0;
      ways_1_metas_101_vld <= 1'b0;
      ways_1_metas_101_tag <= 51'h0;
      ways_1_metas_101_mru <= 1'b0;
      ways_1_metas_102_vld <= 1'b0;
      ways_1_metas_102_tag <= 51'h0;
      ways_1_metas_102_mru <= 1'b0;
      ways_1_metas_103_vld <= 1'b0;
      ways_1_metas_103_tag <= 51'h0;
      ways_1_metas_103_mru <= 1'b0;
      ways_1_metas_104_vld <= 1'b0;
      ways_1_metas_104_tag <= 51'h0;
      ways_1_metas_104_mru <= 1'b0;
      ways_1_metas_105_vld <= 1'b0;
      ways_1_metas_105_tag <= 51'h0;
      ways_1_metas_105_mru <= 1'b0;
      ways_1_metas_106_vld <= 1'b0;
      ways_1_metas_106_tag <= 51'h0;
      ways_1_metas_106_mru <= 1'b0;
      ways_1_metas_107_vld <= 1'b0;
      ways_1_metas_107_tag <= 51'h0;
      ways_1_metas_107_mru <= 1'b0;
      ways_1_metas_108_vld <= 1'b0;
      ways_1_metas_108_tag <= 51'h0;
      ways_1_metas_108_mru <= 1'b0;
      ways_1_metas_109_vld <= 1'b0;
      ways_1_metas_109_tag <= 51'h0;
      ways_1_metas_109_mru <= 1'b0;
      ways_1_metas_110_vld <= 1'b0;
      ways_1_metas_110_tag <= 51'h0;
      ways_1_metas_110_mru <= 1'b0;
      ways_1_metas_111_vld <= 1'b0;
      ways_1_metas_111_tag <= 51'h0;
      ways_1_metas_111_mru <= 1'b0;
      ways_1_metas_112_vld <= 1'b0;
      ways_1_metas_112_tag <= 51'h0;
      ways_1_metas_112_mru <= 1'b0;
      ways_1_metas_113_vld <= 1'b0;
      ways_1_metas_113_tag <= 51'h0;
      ways_1_metas_113_mru <= 1'b0;
      ways_1_metas_114_vld <= 1'b0;
      ways_1_metas_114_tag <= 51'h0;
      ways_1_metas_114_mru <= 1'b0;
      ways_1_metas_115_vld <= 1'b0;
      ways_1_metas_115_tag <= 51'h0;
      ways_1_metas_115_mru <= 1'b0;
      ways_1_metas_116_vld <= 1'b0;
      ways_1_metas_116_tag <= 51'h0;
      ways_1_metas_116_mru <= 1'b0;
      ways_1_metas_117_vld <= 1'b0;
      ways_1_metas_117_tag <= 51'h0;
      ways_1_metas_117_mru <= 1'b0;
      ways_1_metas_118_vld <= 1'b0;
      ways_1_metas_118_tag <= 51'h0;
      ways_1_metas_118_mru <= 1'b0;
      ways_1_metas_119_vld <= 1'b0;
      ways_1_metas_119_tag <= 51'h0;
      ways_1_metas_119_mru <= 1'b0;
      ways_1_metas_120_vld <= 1'b0;
      ways_1_metas_120_tag <= 51'h0;
      ways_1_metas_120_mru <= 1'b0;
      ways_1_metas_121_vld <= 1'b0;
      ways_1_metas_121_tag <= 51'h0;
      ways_1_metas_121_mru <= 1'b0;
      ways_1_metas_122_vld <= 1'b0;
      ways_1_metas_122_tag <= 51'h0;
      ways_1_metas_122_mru <= 1'b0;
      ways_1_metas_123_vld <= 1'b0;
      ways_1_metas_123_tag <= 51'h0;
      ways_1_metas_123_mru <= 1'b0;
      ways_1_metas_124_vld <= 1'b0;
      ways_1_metas_124_tag <= 51'h0;
      ways_1_metas_124_mru <= 1'b0;
      ways_1_metas_125_vld <= 1'b0;
      ways_1_metas_125_tag <= 51'h0;
      ways_1_metas_125_mru <= 1'b0;
      ways_1_metas_126_vld <= 1'b0;
      ways_1_metas_126_tag <= 51'h0;
      ways_1_metas_126_mru <= 1'b0;
      ways_1_metas_127_vld <= 1'b0;
      ways_1_metas_127_tag <= 51'h0;
      ways_1_metas_127_mru <= 1'b0;
      ways_2_metas_0_vld <= 1'b0;
      ways_2_metas_0_tag <= 51'h0;
      ways_2_metas_0_mru <= 1'b0;
      ways_2_metas_1_vld <= 1'b0;
      ways_2_metas_1_tag <= 51'h0;
      ways_2_metas_1_mru <= 1'b0;
      ways_2_metas_2_vld <= 1'b0;
      ways_2_metas_2_tag <= 51'h0;
      ways_2_metas_2_mru <= 1'b0;
      ways_2_metas_3_vld <= 1'b0;
      ways_2_metas_3_tag <= 51'h0;
      ways_2_metas_3_mru <= 1'b0;
      ways_2_metas_4_vld <= 1'b0;
      ways_2_metas_4_tag <= 51'h0;
      ways_2_metas_4_mru <= 1'b0;
      ways_2_metas_5_vld <= 1'b0;
      ways_2_metas_5_tag <= 51'h0;
      ways_2_metas_5_mru <= 1'b0;
      ways_2_metas_6_vld <= 1'b0;
      ways_2_metas_6_tag <= 51'h0;
      ways_2_metas_6_mru <= 1'b0;
      ways_2_metas_7_vld <= 1'b0;
      ways_2_metas_7_tag <= 51'h0;
      ways_2_metas_7_mru <= 1'b0;
      ways_2_metas_8_vld <= 1'b0;
      ways_2_metas_8_tag <= 51'h0;
      ways_2_metas_8_mru <= 1'b0;
      ways_2_metas_9_vld <= 1'b0;
      ways_2_metas_9_tag <= 51'h0;
      ways_2_metas_9_mru <= 1'b0;
      ways_2_metas_10_vld <= 1'b0;
      ways_2_metas_10_tag <= 51'h0;
      ways_2_metas_10_mru <= 1'b0;
      ways_2_metas_11_vld <= 1'b0;
      ways_2_metas_11_tag <= 51'h0;
      ways_2_metas_11_mru <= 1'b0;
      ways_2_metas_12_vld <= 1'b0;
      ways_2_metas_12_tag <= 51'h0;
      ways_2_metas_12_mru <= 1'b0;
      ways_2_metas_13_vld <= 1'b0;
      ways_2_metas_13_tag <= 51'h0;
      ways_2_metas_13_mru <= 1'b0;
      ways_2_metas_14_vld <= 1'b0;
      ways_2_metas_14_tag <= 51'h0;
      ways_2_metas_14_mru <= 1'b0;
      ways_2_metas_15_vld <= 1'b0;
      ways_2_metas_15_tag <= 51'h0;
      ways_2_metas_15_mru <= 1'b0;
      ways_2_metas_16_vld <= 1'b0;
      ways_2_metas_16_tag <= 51'h0;
      ways_2_metas_16_mru <= 1'b0;
      ways_2_metas_17_vld <= 1'b0;
      ways_2_metas_17_tag <= 51'h0;
      ways_2_metas_17_mru <= 1'b0;
      ways_2_metas_18_vld <= 1'b0;
      ways_2_metas_18_tag <= 51'h0;
      ways_2_metas_18_mru <= 1'b0;
      ways_2_metas_19_vld <= 1'b0;
      ways_2_metas_19_tag <= 51'h0;
      ways_2_metas_19_mru <= 1'b0;
      ways_2_metas_20_vld <= 1'b0;
      ways_2_metas_20_tag <= 51'h0;
      ways_2_metas_20_mru <= 1'b0;
      ways_2_metas_21_vld <= 1'b0;
      ways_2_metas_21_tag <= 51'h0;
      ways_2_metas_21_mru <= 1'b0;
      ways_2_metas_22_vld <= 1'b0;
      ways_2_metas_22_tag <= 51'h0;
      ways_2_metas_22_mru <= 1'b0;
      ways_2_metas_23_vld <= 1'b0;
      ways_2_metas_23_tag <= 51'h0;
      ways_2_metas_23_mru <= 1'b0;
      ways_2_metas_24_vld <= 1'b0;
      ways_2_metas_24_tag <= 51'h0;
      ways_2_metas_24_mru <= 1'b0;
      ways_2_metas_25_vld <= 1'b0;
      ways_2_metas_25_tag <= 51'h0;
      ways_2_metas_25_mru <= 1'b0;
      ways_2_metas_26_vld <= 1'b0;
      ways_2_metas_26_tag <= 51'h0;
      ways_2_metas_26_mru <= 1'b0;
      ways_2_metas_27_vld <= 1'b0;
      ways_2_metas_27_tag <= 51'h0;
      ways_2_metas_27_mru <= 1'b0;
      ways_2_metas_28_vld <= 1'b0;
      ways_2_metas_28_tag <= 51'h0;
      ways_2_metas_28_mru <= 1'b0;
      ways_2_metas_29_vld <= 1'b0;
      ways_2_metas_29_tag <= 51'h0;
      ways_2_metas_29_mru <= 1'b0;
      ways_2_metas_30_vld <= 1'b0;
      ways_2_metas_30_tag <= 51'h0;
      ways_2_metas_30_mru <= 1'b0;
      ways_2_metas_31_vld <= 1'b0;
      ways_2_metas_31_tag <= 51'h0;
      ways_2_metas_31_mru <= 1'b0;
      ways_2_metas_32_vld <= 1'b0;
      ways_2_metas_32_tag <= 51'h0;
      ways_2_metas_32_mru <= 1'b0;
      ways_2_metas_33_vld <= 1'b0;
      ways_2_metas_33_tag <= 51'h0;
      ways_2_metas_33_mru <= 1'b0;
      ways_2_metas_34_vld <= 1'b0;
      ways_2_metas_34_tag <= 51'h0;
      ways_2_metas_34_mru <= 1'b0;
      ways_2_metas_35_vld <= 1'b0;
      ways_2_metas_35_tag <= 51'h0;
      ways_2_metas_35_mru <= 1'b0;
      ways_2_metas_36_vld <= 1'b0;
      ways_2_metas_36_tag <= 51'h0;
      ways_2_metas_36_mru <= 1'b0;
      ways_2_metas_37_vld <= 1'b0;
      ways_2_metas_37_tag <= 51'h0;
      ways_2_metas_37_mru <= 1'b0;
      ways_2_metas_38_vld <= 1'b0;
      ways_2_metas_38_tag <= 51'h0;
      ways_2_metas_38_mru <= 1'b0;
      ways_2_metas_39_vld <= 1'b0;
      ways_2_metas_39_tag <= 51'h0;
      ways_2_metas_39_mru <= 1'b0;
      ways_2_metas_40_vld <= 1'b0;
      ways_2_metas_40_tag <= 51'h0;
      ways_2_metas_40_mru <= 1'b0;
      ways_2_metas_41_vld <= 1'b0;
      ways_2_metas_41_tag <= 51'h0;
      ways_2_metas_41_mru <= 1'b0;
      ways_2_metas_42_vld <= 1'b0;
      ways_2_metas_42_tag <= 51'h0;
      ways_2_metas_42_mru <= 1'b0;
      ways_2_metas_43_vld <= 1'b0;
      ways_2_metas_43_tag <= 51'h0;
      ways_2_metas_43_mru <= 1'b0;
      ways_2_metas_44_vld <= 1'b0;
      ways_2_metas_44_tag <= 51'h0;
      ways_2_metas_44_mru <= 1'b0;
      ways_2_metas_45_vld <= 1'b0;
      ways_2_metas_45_tag <= 51'h0;
      ways_2_metas_45_mru <= 1'b0;
      ways_2_metas_46_vld <= 1'b0;
      ways_2_metas_46_tag <= 51'h0;
      ways_2_metas_46_mru <= 1'b0;
      ways_2_metas_47_vld <= 1'b0;
      ways_2_metas_47_tag <= 51'h0;
      ways_2_metas_47_mru <= 1'b0;
      ways_2_metas_48_vld <= 1'b0;
      ways_2_metas_48_tag <= 51'h0;
      ways_2_metas_48_mru <= 1'b0;
      ways_2_metas_49_vld <= 1'b0;
      ways_2_metas_49_tag <= 51'h0;
      ways_2_metas_49_mru <= 1'b0;
      ways_2_metas_50_vld <= 1'b0;
      ways_2_metas_50_tag <= 51'h0;
      ways_2_metas_50_mru <= 1'b0;
      ways_2_metas_51_vld <= 1'b0;
      ways_2_metas_51_tag <= 51'h0;
      ways_2_metas_51_mru <= 1'b0;
      ways_2_metas_52_vld <= 1'b0;
      ways_2_metas_52_tag <= 51'h0;
      ways_2_metas_52_mru <= 1'b0;
      ways_2_metas_53_vld <= 1'b0;
      ways_2_metas_53_tag <= 51'h0;
      ways_2_metas_53_mru <= 1'b0;
      ways_2_metas_54_vld <= 1'b0;
      ways_2_metas_54_tag <= 51'h0;
      ways_2_metas_54_mru <= 1'b0;
      ways_2_metas_55_vld <= 1'b0;
      ways_2_metas_55_tag <= 51'h0;
      ways_2_metas_55_mru <= 1'b0;
      ways_2_metas_56_vld <= 1'b0;
      ways_2_metas_56_tag <= 51'h0;
      ways_2_metas_56_mru <= 1'b0;
      ways_2_metas_57_vld <= 1'b0;
      ways_2_metas_57_tag <= 51'h0;
      ways_2_metas_57_mru <= 1'b0;
      ways_2_metas_58_vld <= 1'b0;
      ways_2_metas_58_tag <= 51'h0;
      ways_2_metas_58_mru <= 1'b0;
      ways_2_metas_59_vld <= 1'b0;
      ways_2_metas_59_tag <= 51'h0;
      ways_2_metas_59_mru <= 1'b0;
      ways_2_metas_60_vld <= 1'b0;
      ways_2_metas_60_tag <= 51'h0;
      ways_2_metas_60_mru <= 1'b0;
      ways_2_metas_61_vld <= 1'b0;
      ways_2_metas_61_tag <= 51'h0;
      ways_2_metas_61_mru <= 1'b0;
      ways_2_metas_62_vld <= 1'b0;
      ways_2_metas_62_tag <= 51'h0;
      ways_2_metas_62_mru <= 1'b0;
      ways_2_metas_63_vld <= 1'b0;
      ways_2_metas_63_tag <= 51'h0;
      ways_2_metas_63_mru <= 1'b0;
      ways_2_metas_64_vld <= 1'b0;
      ways_2_metas_64_tag <= 51'h0;
      ways_2_metas_64_mru <= 1'b0;
      ways_2_metas_65_vld <= 1'b0;
      ways_2_metas_65_tag <= 51'h0;
      ways_2_metas_65_mru <= 1'b0;
      ways_2_metas_66_vld <= 1'b0;
      ways_2_metas_66_tag <= 51'h0;
      ways_2_metas_66_mru <= 1'b0;
      ways_2_metas_67_vld <= 1'b0;
      ways_2_metas_67_tag <= 51'h0;
      ways_2_metas_67_mru <= 1'b0;
      ways_2_metas_68_vld <= 1'b0;
      ways_2_metas_68_tag <= 51'h0;
      ways_2_metas_68_mru <= 1'b0;
      ways_2_metas_69_vld <= 1'b0;
      ways_2_metas_69_tag <= 51'h0;
      ways_2_metas_69_mru <= 1'b0;
      ways_2_metas_70_vld <= 1'b0;
      ways_2_metas_70_tag <= 51'h0;
      ways_2_metas_70_mru <= 1'b0;
      ways_2_metas_71_vld <= 1'b0;
      ways_2_metas_71_tag <= 51'h0;
      ways_2_metas_71_mru <= 1'b0;
      ways_2_metas_72_vld <= 1'b0;
      ways_2_metas_72_tag <= 51'h0;
      ways_2_metas_72_mru <= 1'b0;
      ways_2_metas_73_vld <= 1'b0;
      ways_2_metas_73_tag <= 51'h0;
      ways_2_metas_73_mru <= 1'b0;
      ways_2_metas_74_vld <= 1'b0;
      ways_2_metas_74_tag <= 51'h0;
      ways_2_metas_74_mru <= 1'b0;
      ways_2_metas_75_vld <= 1'b0;
      ways_2_metas_75_tag <= 51'h0;
      ways_2_metas_75_mru <= 1'b0;
      ways_2_metas_76_vld <= 1'b0;
      ways_2_metas_76_tag <= 51'h0;
      ways_2_metas_76_mru <= 1'b0;
      ways_2_metas_77_vld <= 1'b0;
      ways_2_metas_77_tag <= 51'h0;
      ways_2_metas_77_mru <= 1'b0;
      ways_2_metas_78_vld <= 1'b0;
      ways_2_metas_78_tag <= 51'h0;
      ways_2_metas_78_mru <= 1'b0;
      ways_2_metas_79_vld <= 1'b0;
      ways_2_metas_79_tag <= 51'h0;
      ways_2_metas_79_mru <= 1'b0;
      ways_2_metas_80_vld <= 1'b0;
      ways_2_metas_80_tag <= 51'h0;
      ways_2_metas_80_mru <= 1'b0;
      ways_2_metas_81_vld <= 1'b0;
      ways_2_metas_81_tag <= 51'h0;
      ways_2_metas_81_mru <= 1'b0;
      ways_2_metas_82_vld <= 1'b0;
      ways_2_metas_82_tag <= 51'h0;
      ways_2_metas_82_mru <= 1'b0;
      ways_2_metas_83_vld <= 1'b0;
      ways_2_metas_83_tag <= 51'h0;
      ways_2_metas_83_mru <= 1'b0;
      ways_2_metas_84_vld <= 1'b0;
      ways_2_metas_84_tag <= 51'h0;
      ways_2_metas_84_mru <= 1'b0;
      ways_2_metas_85_vld <= 1'b0;
      ways_2_metas_85_tag <= 51'h0;
      ways_2_metas_85_mru <= 1'b0;
      ways_2_metas_86_vld <= 1'b0;
      ways_2_metas_86_tag <= 51'h0;
      ways_2_metas_86_mru <= 1'b0;
      ways_2_metas_87_vld <= 1'b0;
      ways_2_metas_87_tag <= 51'h0;
      ways_2_metas_87_mru <= 1'b0;
      ways_2_metas_88_vld <= 1'b0;
      ways_2_metas_88_tag <= 51'h0;
      ways_2_metas_88_mru <= 1'b0;
      ways_2_metas_89_vld <= 1'b0;
      ways_2_metas_89_tag <= 51'h0;
      ways_2_metas_89_mru <= 1'b0;
      ways_2_metas_90_vld <= 1'b0;
      ways_2_metas_90_tag <= 51'h0;
      ways_2_metas_90_mru <= 1'b0;
      ways_2_metas_91_vld <= 1'b0;
      ways_2_metas_91_tag <= 51'h0;
      ways_2_metas_91_mru <= 1'b0;
      ways_2_metas_92_vld <= 1'b0;
      ways_2_metas_92_tag <= 51'h0;
      ways_2_metas_92_mru <= 1'b0;
      ways_2_metas_93_vld <= 1'b0;
      ways_2_metas_93_tag <= 51'h0;
      ways_2_metas_93_mru <= 1'b0;
      ways_2_metas_94_vld <= 1'b0;
      ways_2_metas_94_tag <= 51'h0;
      ways_2_metas_94_mru <= 1'b0;
      ways_2_metas_95_vld <= 1'b0;
      ways_2_metas_95_tag <= 51'h0;
      ways_2_metas_95_mru <= 1'b0;
      ways_2_metas_96_vld <= 1'b0;
      ways_2_metas_96_tag <= 51'h0;
      ways_2_metas_96_mru <= 1'b0;
      ways_2_metas_97_vld <= 1'b0;
      ways_2_metas_97_tag <= 51'h0;
      ways_2_metas_97_mru <= 1'b0;
      ways_2_metas_98_vld <= 1'b0;
      ways_2_metas_98_tag <= 51'h0;
      ways_2_metas_98_mru <= 1'b0;
      ways_2_metas_99_vld <= 1'b0;
      ways_2_metas_99_tag <= 51'h0;
      ways_2_metas_99_mru <= 1'b0;
      ways_2_metas_100_vld <= 1'b0;
      ways_2_metas_100_tag <= 51'h0;
      ways_2_metas_100_mru <= 1'b0;
      ways_2_metas_101_vld <= 1'b0;
      ways_2_metas_101_tag <= 51'h0;
      ways_2_metas_101_mru <= 1'b0;
      ways_2_metas_102_vld <= 1'b0;
      ways_2_metas_102_tag <= 51'h0;
      ways_2_metas_102_mru <= 1'b0;
      ways_2_metas_103_vld <= 1'b0;
      ways_2_metas_103_tag <= 51'h0;
      ways_2_metas_103_mru <= 1'b0;
      ways_2_metas_104_vld <= 1'b0;
      ways_2_metas_104_tag <= 51'h0;
      ways_2_metas_104_mru <= 1'b0;
      ways_2_metas_105_vld <= 1'b0;
      ways_2_metas_105_tag <= 51'h0;
      ways_2_metas_105_mru <= 1'b0;
      ways_2_metas_106_vld <= 1'b0;
      ways_2_metas_106_tag <= 51'h0;
      ways_2_metas_106_mru <= 1'b0;
      ways_2_metas_107_vld <= 1'b0;
      ways_2_metas_107_tag <= 51'h0;
      ways_2_metas_107_mru <= 1'b0;
      ways_2_metas_108_vld <= 1'b0;
      ways_2_metas_108_tag <= 51'h0;
      ways_2_metas_108_mru <= 1'b0;
      ways_2_metas_109_vld <= 1'b0;
      ways_2_metas_109_tag <= 51'h0;
      ways_2_metas_109_mru <= 1'b0;
      ways_2_metas_110_vld <= 1'b0;
      ways_2_metas_110_tag <= 51'h0;
      ways_2_metas_110_mru <= 1'b0;
      ways_2_metas_111_vld <= 1'b0;
      ways_2_metas_111_tag <= 51'h0;
      ways_2_metas_111_mru <= 1'b0;
      ways_2_metas_112_vld <= 1'b0;
      ways_2_metas_112_tag <= 51'h0;
      ways_2_metas_112_mru <= 1'b0;
      ways_2_metas_113_vld <= 1'b0;
      ways_2_metas_113_tag <= 51'h0;
      ways_2_metas_113_mru <= 1'b0;
      ways_2_metas_114_vld <= 1'b0;
      ways_2_metas_114_tag <= 51'h0;
      ways_2_metas_114_mru <= 1'b0;
      ways_2_metas_115_vld <= 1'b0;
      ways_2_metas_115_tag <= 51'h0;
      ways_2_metas_115_mru <= 1'b0;
      ways_2_metas_116_vld <= 1'b0;
      ways_2_metas_116_tag <= 51'h0;
      ways_2_metas_116_mru <= 1'b0;
      ways_2_metas_117_vld <= 1'b0;
      ways_2_metas_117_tag <= 51'h0;
      ways_2_metas_117_mru <= 1'b0;
      ways_2_metas_118_vld <= 1'b0;
      ways_2_metas_118_tag <= 51'h0;
      ways_2_metas_118_mru <= 1'b0;
      ways_2_metas_119_vld <= 1'b0;
      ways_2_metas_119_tag <= 51'h0;
      ways_2_metas_119_mru <= 1'b0;
      ways_2_metas_120_vld <= 1'b0;
      ways_2_metas_120_tag <= 51'h0;
      ways_2_metas_120_mru <= 1'b0;
      ways_2_metas_121_vld <= 1'b0;
      ways_2_metas_121_tag <= 51'h0;
      ways_2_metas_121_mru <= 1'b0;
      ways_2_metas_122_vld <= 1'b0;
      ways_2_metas_122_tag <= 51'h0;
      ways_2_metas_122_mru <= 1'b0;
      ways_2_metas_123_vld <= 1'b0;
      ways_2_metas_123_tag <= 51'h0;
      ways_2_metas_123_mru <= 1'b0;
      ways_2_metas_124_vld <= 1'b0;
      ways_2_metas_124_tag <= 51'h0;
      ways_2_metas_124_mru <= 1'b0;
      ways_2_metas_125_vld <= 1'b0;
      ways_2_metas_125_tag <= 51'h0;
      ways_2_metas_125_mru <= 1'b0;
      ways_2_metas_126_vld <= 1'b0;
      ways_2_metas_126_tag <= 51'h0;
      ways_2_metas_126_mru <= 1'b0;
      ways_2_metas_127_vld <= 1'b0;
      ways_2_metas_127_tag <= 51'h0;
      ways_2_metas_127_mru <= 1'b0;
      ways_3_metas_0_vld <= 1'b0;
      ways_3_metas_0_tag <= 51'h0;
      ways_3_metas_0_mru <= 1'b0;
      ways_3_metas_1_vld <= 1'b0;
      ways_3_metas_1_tag <= 51'h0;
      ways_3_metas_1_mru <= 1'b0;
      ways_3_metas_2_vld <= 1'b0;
      ways_3_metas_2_tag <= 51'h0;
      ways_3_metas_2_mru <= 1'b0;
      ways_3_metas_3_vld <= 1'b0;
      ways_3_metas_3_tag <= 51'h0;
      ways_3_metas_3_mru <= 1'b0;
      ways_3_metas_4_vld <= 1'b0;
      ways_3_metas_4_tag <= 51'h0;
      ways_3_metas_4_mru <= 1'b0;
      ways_3_metas_5_vld <= 1'b0;
      ways_3_metas_5_tag <= 51'h0;
      ways_3_metas_5_mru <= 1'b0;
      ways_3_metas_6_vld <= 1'b0;
      ways_3_metas_6_tag <= 51'h0;
      ways_3_metas_6_mru <= 1'b0;
      ways_3_metas_7_vld <= 1'b0;
      ways_3_metas_7_tag <= 51'h0;
      ways_3_metas_7_mru <= 1'b0;
      ways_3_metas_8_vld <= 1'b0;
      ways_3_metas_8_tag <= 51'h0;
      ways_3_metas_8_mru <= 1'b0;
      ways_3_metas_9_vld <= 1'b0;
      ways_3_metas_9_tag <= 51'h0;
      ways_3_metas_9_mru <= 1'b0;
      ways_3_metas_10_vld <= 1'b0;
      ways_3_metas_10_tag <= 51'h0;
      ways_3_metas_10_mru <= 1'b0;
      ways_3_metas_11_vld <= 1'b0;
      ways_3_metas_11_tag <= 51'h0;
      ways_3_metas_11_mru <= 1'b0;
      ways_3_metas_12_vld <= 1'b0;
      ways_3_metas_12_tag <= 51'h0;
      ways_3_metas_12_mru <= 1'b0;
      ways_3_metas_13_vld <= 1'b0;
      ways_3_metas_13_tag <= 51'h0;
      ways_3_metas_13_mru <= 1'b0;
      ways_3_metas_14_vld <= 1'b0;
      ways_3_metas_14_tag <= 51'h0;
      ways_3_metas_14_mru <= 1'b0;
      ways_3_metas_15_vld <= 1'b0;
      ways_3_metas_15_tag <= 51'h0;
      ways_3_metas_15_mru <= 1'b0;
      ways_3_metas_16_vld <= 1'b0;
      ways_3_metas_16_tag <= 51'h0;
      ways_3_metas_16_mru <= 1'b0;
      ways_3_metas_17_vld <= 1'b0;
      ways_3_metas_17_tag <= 51'h0;
      ways_3_metas_17_mru <= 1'b0;
      ways_3_metas_18_vld <= 1'b0;
      ways_3_metas_18_tag <= 51'h0;
      ways_3_metas_18_mru <= 1'b0;
      ways_3_metas_19_vld <= 1'b0;
      ways_3_metas_19_tag <= 51'h0;
      ways_3_metas_19_mru <= 1'b0;
      ways_3_metas_20_vld <= 1'b0;
      ways_3_metas_20_tag <= 51'h0;
      ways_3_metas_20_mru <= 1'b0;
      ways_3_metas_21_vld <= 1'b0;
      ways_3_metas_21_tag <= 51'h0;
      ways_3_metas_21_mru <= 1'b0;
      ways_3_metas_22_vld <= 1'b0;
      ways_3_metas_22_tag <= 51'h0;
      ways_3_metas_22_mru <= 1'b0;
      ways_3_metas_23_vld <= 1'b0;
      ways_3_metas_23_tag <= 51'h0;
      ways_3_metas_23_mru <= 1'b0;
      ways_3_metas_24_vld <= 1'b0;
      ways_3_metas_24_tag <= 51'h0;
      ways_3_metas_24_mru <= 1'b0;
      ways_3_metas_25_vld <= 1'b0;
      ways_3_metas_25_tag <= 51'h0;
      ways_3_metas_25_mru <= 1'b0;
      ways_3_metas_26_vld <= 1'b0;
      ways_3_metas_26_tag <= 51'h0;
      ways_3_metas_26_mru <= 1'b0;
      ways_3_metas_27_vld <= 1'b0;
      ways_3_metas_27_tag <= 51'h0;
      ways_3_metas_27_mru <= 1'b0;
      ways_3_metas_28_vld <= 1'b0;
      ways_3_metas_28_tag <= 51'h0;
      ways_3_metas_28_mru <= 1'b0;
      ways_3_metas_29_vld <= 1'b0;
      ways_3_metas_29_tag <= 51'h0;
      ways_3_metas_29_mru <= 1'b0;
      ways_3_metas_30_vld <= 1'b0;
      ways_3_metas_30_tag <= 51'h0;
      ways_3_metas_30_mru <= 1'b0;
      ways_3_metas_31_vld <= 1'b0;
      ways_3_metas_31_tag <= 51'h0;
      ways_3_metas_31_mru <= 1'b0;
      ways_3_metas_32_vld <= 1'b0;
      ways_3_metas_32_tag <= 51'h0;
      ways_3_metas_32_mru <= 1'b0;
      ways_3_metas_33_vld <= 1'b0;
      ways_3_metas_33_tag <= 51'h0;
      ways_3_metas_33_mru <= 1'b0;
      ways_3_metas_34_vld <= 1'b0;
      ways_3_metas_34_tag <= 51'h0;
      ways_3_metas_34_mru <= 1'b0;
      ways_3_metas_35_vld <= 1'b0;
      ways_3_metas_35_tag <= 51'h0;
      ways_3_metas_35_mru <= 1'b0;
      ways_3_metas_36_vld <= 1'b0;
      ways_3_metas_36_tag <= 51'h0;
      ways_3_metas_36_mru <= 1'b0;
      ways_3_metas_37_vld <= 1'b0;
      ways_3_metas_37_tag <= 51'h0;
      ways_3_metas_37_mru <= 1'b0;
      ways_3_metas_38_vld <= 1'b0;
      ways_3_metas_38_tag <= 51'h0;
      ways_3_metas_38_mru <= 1'b0;
      ways_3_metas_39_vld <= 1'b0;
      ways_3_metas_39_tag <= 51'h0;
      ways_3_metas_39_mru <= 1'b0;
      ways_3_metas_40_vld <= 1'b0;
      ways_3_metas_40_tag <= 51'h0;
      ways_3_metas_40_mru <= 1'b0;
      ways_3_metas_41_vld <= 1'b0;
      ways_3_metas_41_tag <= 51'h0;
      ways_3_metas_41_mru <= 1'b0;
      ways_3_metas_42_vld <= 1'b0;
      ways_3_metas_42_tag <= 51'h0;
      ways_3_metas_42_mru <= 1'b0;
      ways_3_metas_43_vld <= 1'b0;
      ways_3_metas_43_tag <= 51'h0;
      ways_3_metas_43_mru <= 1'b0;
      ways_3_metas_44_vld <= 1'b0;
      ways_3_metas_44_tag <= 51'h0;
      ways_3_metas_44_mru <= 1'b0;
      ways_3_metas_45_vld <= 1'b0;
      ways_3_metas_45_tag <= 51'h0;
      ways_3_metas_45_mru <= 1'b0;
      ways_3_metas_46_vld <= 1'b0;
      ways_3_metas_46_tag <= 51'h0;
      ways_3_metas_46_mru <= 1'b0;
      ways_3_metas_47_vld <= 1'b0;
      ways_3_metas_47_tag <= 51'h0;
      ways_3_metas_47_mru <= 1'b0;
      ways_3_metas_48_vld <= 1'b0;
      ways_3_metas_48_tag <= 51'h0;
      ways_3_metas_48_mru <= 1'b0;
      ways_3_metas_49_vld <= 1'b0;
      ways_3_metas_49_tag <= 51'h0;
      ways_3_metas_49_mru <= 1'b0;
      ways_3_metas_50_vld <= 1'b0;
      ways_3_metas_50_tag <= 51'h0;
      ways_3_metas_50_mru <= 1'b0;
      ways_3_metas_51_vld <= 1'b0;
      ways_3_metas_51_tag <= 51'h0;
      ways_3_metas_51_mru <= 1'b0;
      ways_3_metas_52_vld <= 1'b0;
      ways_3_metas_52_tag <= 51'h0;
      ways_3_metas_52_mru <= 1'b0;
      ways_3_metas_53_vld <= 1'b0;
      ways_3_metas_53_tag <= 51'h0;
      ways_3_metas_53_mru <= 1'b0;
      ways_3_metas_54_vld <= 1'b0;
      ways_3_metas_54_tag <= 51'h0;
      ways_3_metas_54_mru <= 1'b0;
      ways_3_metas_55_vld <= 1'b0;
      ways_3_metas_55_tag <= 51'h0;
      ways_3_metas_55_mru <= 1'b0;
      ways_3_metas_56_vld <= 1'b0;
      ways_3_metas_56_tag <= 51'h0;
      ways_3_metas_56_mru <= 1'b0;
      ways_3_metas_57_vld <= 1'b0;
      ways_3_metas_57_tag <= 51'h0;
      ways_3_metas_57_mru <= 1'b0;
      ways_3_metas_58_vld <= 1'b0;
      ways_3_metas_58_tag <= 51'h0;
      ways_3_metas_58_mru <= 1'b0;
      ways_3_metas_59_vld <= 1'b0;
      ways_3_metas_59_tag <= 51'h0;
      ways_3_metas_59_mru <= 1'b0;
      ways_3_metas_60_vld <= 1'b0;
      ways_3_metas_60_tag <= 51'h0;
      ways_3_metas_60_mru <= 1'b0;
      ways_3_metas_61_vld <= 1'b0;
      ways_3_metas_61_tag <= 51'h0;
      ways_3_metas_61_mru <= 1'b0;
      ways_3_metas_62_vld <= 1'b0;
      ways_3_metas_62_tag <= 51'h0;
      ways_3_metas_62_mru <= 1'b0;
      ways_3_metas_63_vld <= 1'b0;
      ways_3_metas_63_tag <= 51'h0;
      ways_3_metas_63_mru <= 1'b0;
      ways_3_metas_64_vld <= 1'b0;
      ways_3_metas_64_tag <= 51'h0;
      ways_3_metas_64_mru <= 1'b0;
      ways_3_metas_65_vld <= 1'b0;
      ways_3_metas_65_tag <= 51'h0;
      ways_3_metas_65_mru <= 1'b0;
      ways_3_metas_66_vld <= 1'b0;
      ways_3_metas_66_tag <= 51'h0;
      ways_3_metas_66_mru <= 1'b0;
      ways_3_metas_67_vld <= 1'b0;
      ways_3_metas_67_tag <= 51'h0;
      ways_3_metas_67_mru <= 1'b0;
      ways_3_metas_68_vld <= 1'b0;
      ways_3_metas_68_tag <= 51'h0;
      ways_3_metas_68_mru <= 1'b0;
      ways_3_metas_69_vld <= 1'b0;
      ways_3_metas_69_tag <= 51'h0;
      ways_3_metas_69_mru <= 1'b0;
      ways_3_metas_70_vld <= 1'b0;
      ways_3_metas_70_tag <= 51'h0;
      ways_3_metas_70_mru <= 1'b0;
      ways_3_metas_71_vld <= 1'b0;
      ways_3_metas_71_tag <= 51'h0;
      ways_3_metas_71_mru <= 1'b0;
      ways_3_metas_72_vld <= 1'b0;
      ways_3_metas_72_tag <= 51'h0;
      ways_3_metas_72_mru <= 1'b0;
      ways_3_metas_73_vld <= 1'b0;
      ways_3_metas_73_tag <= 51'h0;
      ways_3_metas_73_mru <= 1'b0;
      ways_3_metas_74_vld <= 1'b0;
      ways_3_metas_74_tag <= 51'h0;
      ways_3_metas_74_mru <= 1'b0;
      ways_3_metas_75_vld <= 1'b0;
      ways_3_metas_75_tag <= 51'h0;
      ways_3_metas_75_mru <= 1'b0;
      ways_3_metas_76_vld <= 1'b0;
      ways_3_metas_76_tag <= 51'h0;
      ways_3_metas_76_mru <= 1'b0;
      ways_3_metas_77_vld <= 1'b0;
      ways_3_metas_77_tag <= 51'h0;
      ways_3_metas_77_mru <= 1'b0;
      ways_3_metas_78_vld <= 1'b0;
      ways_3_metas_78_tag <= 51'h0;
      ways_3_metas_78_mru <= 1'b0;
      ways_3_metas_79_vld <= 1'b0;
      ways_3_metas_79_tag <= 51'h0;
      ways_3_metas_79_mru <= 1'b0;
      ways_3_metas_80_vld <= 1'b0;
      ways_3_metas_80_tag <= 51'h0;
      ways_3_metas_80_mru <= 1'b0;
      ways_3_metas_81_vld <= 1'b0;
      ways_3_metas_81_tag <= 51'h0;
      ways_3_metas_81_mru <= 1'b0;
      ways_3_metas_82_vld <= 1'b0;
      ways_3_metas_82_tag <= 51'h0;
      ways_3_metas_82_mru <= 1'b0;
      ways_3_metas_83_vld <= 1'b0;
      ways_3_metas_83_tag <= 51'h0;
      ways_3_metas_83_mru <= 1'b0;
      ways_3_metas_84_vld <= 1'b0;
      ways_3_metas_84_tag <= 51'h0;
      ways_3_metas_84_mru <= 1'b0;
      ways_3_metas_85_vld <= 1'b0;
      ways_3_metas_85_tag <= 51'h0;
      ways_3_metas_85_mru <= 1'b0;
      ways_3_metas_86_vld <= 1'b0;
      ways_3_metas_86_tag <= 51'h0;
      ways_3_metas_86_mru <= 1'b0;
      ways_3_metas_87_vld <= 1'b0;
      ways_3_metas_87_tag <= 51'h0;
      ways_3_metas_87_mru <= 1'b0;
      ways_3_metas_88_vld <= 1'b0;
      ways_3_metas_88_tag <= 51'h0;
      ways_3_metas_88_mru <= 1'b0;
      ways_3_metas_89_vld <= 1'b0;
      ways_3_metas_89_tag <= 51'h0;
      ways_3_metas_89_mru <= 1'b0;
      ways_3_metas_90_vld <= 1'b0;
      ways_3_metas_90_tag <= 51'h0;
      ways_3_metas_90_mru <= 1'b0;
      ways_3_metas_91_vld <= 1'b0;
      ways_3_metas_91_tag <= 51'h0;
      ways_3_metas_91_mru <= 1'b0;
      ways_3_metas_92_vld <= 1'b0;
      ways_3_metas_92_tag <= 51'h0;
      ways_3_metas_92_mru <= 1'b0;
      ways_3_metas_93_vld <= 1'b0;
      ways_3_metas_93_tag <= 51'h0;
      ways_3_metas_93_mru <= 1'b0;
      ways_3_metas_94_vld <= 1'b0;
      ways_3_metas_94_tag <= 51'h0;
      ways_3_metas_94_mru <= 1'b0;
      ways_3_metas_95_vld <= 1'b0;
      ways_3_metas_95_tag <= 51'h0;
      ways_3_metas_95_mru <= 1'b0;
      ways_3_metas_96_vld <= 1'b0;
      ways_3_metas_96_tag <= 51'h0;
      ways_3_metas_96_mru <= 1'b0;
      ways_3_metas_97_vld <= 1'b0;
      ways_3_metas_97_tag <= 51'h0;
      ways_3_metas_97_mru <= 1'b0;
      ways_3_metas_98_vld <= 1'b0;
      ways_3_metas_98_tag <= 51'h0;
      ways_3_metas_98_mru <= 1'b0;
      ways_3_metas_99_vld <= 1'b0;
      ways_3_metas_99_tag <= 51'h0;
      ways_3_metas_99_mru <= 1'b0;
      ways_3_metas_100_vld <= 1'b0;
      ways_3_metas_100_tag <= 51'h0;
      ways_3_metas_100_mru <= 1'b0;
      ways_3_metas_101_vld <= 1'b0;
      ways_3_metas_101_tag <= 51'h0;
      ways_3_metas_101_mru <= 1'b0;
      ways_3_metas_102_vld <= 1'b0;
      ways_3_metas_102_tag <= 51'h0;
      ways_3_metas_102_mru <= 1'b0;
      ways_3_metas_103_vld <= 1'b0;
      ways_3_metas_103_tag <= 51'h0;
      ways_3_metas_103_mru <= 1'b0;
      ways_3_metas_104_vld <= 1'b0;
      ways_3_metas_104_tag <= 51'h0;
      ways_3_metas_104_mru <= 1'b0;
      ways_3_metas_105_vld <= 1'b0;
      ways_3_metas_105_tag <= 51'h0;
      ways_3_metas_105_mru <= 1'b0;
      ways_3_metas_106_vld <= 1'b0;
      ways_3_metas_106_tag <= 51'h0;
      ways_3_metas_106_mru <= 1'b0;
      ways_3_metas_107_vld <= 1'b0;
      ways_3_metas_107_tag <= 51'h0;
      ways_3_metas_107_mru <= 1'b0;
      ways_3_metas_108_vld <= 1'b0;
      ways_3_metas_108_tag <= 51'h0;
      ways_3_metas_108_mru <= 1'b0;
      ways_3_metas_109_vld <= 1'b0;
      ways_3_metas_109_tag <= 51'h0;
      ways_3_metas_109_mru <= 1'b0;
      ways_3_metas_110_vld <= 1'b0;
      ways_3_metas_110_tag <= 51'h0;
      ways_3_metas_110_mru <= 1'b0;
      ways_3_metas_111_vld <= 1'b0;
      ways_3_metas_111_tag <= 51'h0;
      ways_3_metas_111_mru <= 1'b0;
      ways_3_metas_112_vld <= 1'b0;
      ways_3_metas_112_tag <= 51'h0;
      ways_3_metas_112_mru <= 1'b0;
      ways_3_metas_113_vld <= 1'b0;
      ways_3_metas_113_tag <= 51'h0;
      ways_3_metas_113_mru <= 1'b0;
      ways_3_metas_114_vld <= 1'b0;
      ways_3_metas_114_tag <= 51'h0;
      ways_3_metas_114_mru <= 1'b0;
      ways_3_metas_115_vld <= 1'b0;
      ways_3_metas_115_tag <= 51'h0;
      ways_3_metas_115_mru <= 1'b0;
      ways_3_metas_116_vld <= 1'b0;
      ways_3_metas_116_tag <= 51'h0;
      ways_3_metas_116_mru <= 1'b0;
      ways_3_metas_117_vld <= 1'b0;
      ways_3_metas_117_tag <= 51'h0;
      ways_3_metas_117_mru <= 1'b0;
      ways_3_metas_118_vld <= 1'b0;
      ways_3_metas_118_tag <= 51'h0;
      ways_3_metas_118_mru <= 1'b0;
      ways_3_metas_119_vld <= 1'b0;
      ways_3_metas_119_tag <= 51'h0;
      ways_3_metas_119_mru <= 1'b0;
      ways_3_metas_120_vld <= 1'b0;
      ways_3_metas_120_tag <= 51'h0;
      ways_3_metas_120_mru <= 1'b0;
      ways_3_metas_121_vld <= 1'b0;
      ways_3_metas_121_tag <= 51'h0;
      ways_3_metas_121_mru <= 1'b0;
      ways_3_metas_122_vld <= 1'b0;
      ways_3_metas_122_tag <= 51'h0;
      ways_3_metas_122_mru <= 1'b0;
      ways_3_metas_123_vld <= 1'b0;
      ways_3_metas_123_tag <= 51'h0;
      ways_3_metas_123_mru <= 1'b0;
      ways_3_metas_124_vld <= 1'b0;
      ways_3_metas_124_tag <= 51'h0;
      ways_3_metas_124_mru <= 1'b0;
      ways_3_metas_125_vld <= 1'b0;
      ways_3_metas_125_tag <= 51'h0;
      ways_3_metas_125_mru <= 1'b0;
      ways_3_metas_126_vld <= 1'b0;
      ways_3_metas_126_tag <= 51'h0;
      ways_3_metas_126_mru <= 1'b0;
      ways_3_metas_127_vld <= 1'b0;
      ways_3_metas_127_tag <= 51'h0;
      ways_3_metas_127_mru <= 1'b0;
      flush_busy <= 1'b0;
      flush_cnt_value <= 7'h0;
      cpu_addr_d1 <= 64'h0;
      cpu_cmd_ready_1 <= 1'b1;
      next_level_cmd_valid_1 <= 1'b0;
      next_level_data_cnt_value <= 3'b000;
    end else begin
      flush_cnt_value <= flush_cnt_valueNext;
      if(cpu_cmd_fire_2) begin
        cpu_addr_d1 <= cpu_cmd_payload_addr;
      end
      next_level_data_cnt_value <= next_level_data_cnt_valueNext;
      if(is_miss) begin
        next_level_cmd_valid_1 <= 1'b1;
      end else begin
        if(next_level_cmd_fire) begin
          next_level_cmd_valid_1 <= 1'b0;
        end
      end
      if(flush) begin
        flush_busy <= 1'b1;
      end else begin
        if(flush_done) begin
          flush_busy <= 1'b0;
        end
      end
      if(flush_busy) begin
        if(_zz_260) begin
          ways_0_metas_0_mru <= 1'b0;
        end
        if(_zz_261) begin
          ways_0_metas_1_mru <= 1'b0;
        end
        if(_zz_262) begin
          ways_0_metas_2_mru <= 1'b0;
        end
        if(_zz_263) begin
          ways_0_metas_3_mru <= 1'b0;
        end
        if(_zz_264) begin
          ways_0_metas_4_mru <= 1'b0;
        end
        if(_zz_265) begin
          ways_0_metas_5_mru <= 1'b0;
        end
        if(_zz_266) begin
          ways_0_metas_6_mru <= 1'b0;
        end
        if(_zz_267) begin
          ways_0_metas_7_mru <= 1'b0;
        end
        if(_zz_268) begin
          ways_0_metas_8_mru <= 1'b0;
        end
        if(_zz_269) begin
          ways_0_metas_9_mru <= 1'b0;
        end
        if(_zz_270) begin
          ways_0_metas_10_mru <= 1'b0;
        end
        if(_zz_271) begin
          ways_0_metas_11_mru <= 1'b0;
        end
        if(_zz_272) begin
          ways_0_metas_12_mru <= 1'b0;
        end
        if(_zz_273) begin
          ways_0_metas_13_mru <= 1'b0;
        end
        if(_zz_274) begin
          ways_0_metas_14_mru <= 1'b0;
        end
        if(_zz_275) begin
          ways_0_metas_15_mru <= 1'b0;
        end
        if(_zz_276) begin
          ways_0_metas_16_mru <= 1'b0;
        end
        if(_zz_277) begin
          ways_0_metas_17_mru <= 1'b0;
        end
        if(_zz_278) begin
          ways_0_metas_18_mru <= 1'b0;
        end
        if(_zz_279) begin
          ways_0_metas_19_mru <= 1'b0;
        end
        if(_zz_280) begin
          ways_0_metas_20_mru <= 1'b0;
        end
        if(_zz_281) begin
          ways_0_metas_21_mru <= 1'b0;
        end
        if(_zz_282) begin
          ways_0_metas_22_mru <= 1'b0;
        end
        if(_zz_283) begin
          ways_0_metas_23_mru <= 1'b0;
        end
        if(_zz_284) begin
          ways_0_metas_24_mru <= 1'b0;
        end
        if(_zz_285) begin
          ways_0_metas_25_mru <= 1'b0;
        end
        if(_zz_286) begin
          ways_0_metas_26_mru <= 1'b0;
        end
        if(_zz_287) begin
          ways_0_metas_27_mru <= 1'b0;
        end
        if(_zz_288) begin
          ways_0_metas_28_mru <= 1'b0;
        end
        if(_zz_289) begin
          ways_0_metas_29_mru <= 1'b0;
        end
        if(_zz_290) begin
          ways_0_metas_30_mru <= 1'b0;
        end
        if(_zz_291) begin
          ways_0_metas_31_mru <= 1'b0;
        end
        if(_zz_292) begin
          ways_0_metas_32_mru <= 1'b0;
        end
        if(_zz_293) begin
          ways_0_metas_33_mru <= 1'b0;
        end
        if(_zz_294) begin
          ways_0_metas_34_mru <= 1'b0;
        end
        if(_zz_295) begin
          ways_0_metas_35_mru <= 1'b0;
        end
        if(_zz_296) begin
          ways_0_metas_36_mru <= 1'b0;
        end
        if(_zz_297) begin
          ways_0_metas_37_mru <= 1'b0;
        end
        if(_zz_298) begin
          ways_0_metas_38_mru <= 1'b0;
        end
        if(_zz_299) begin
          ways_0_metas_39_mru <= 1'b0;
        end
        if(_zz_300) begin
          ways_0_metas_40_mru <= 1'b0;
        end
        if(_zz_301) begin
          ways_0_metas_41_mru <= 1'b0;
        end
        if(_zz_302) begin
          ways_0_metas_42_mru <= 1'b0;
        end
        if(_zz_303) begin
          ways_0_metas_43_mru <= 1'b0;
        end
        if(_zz_304) begin
          ways_0_metas_44_mru <= 1'b0;
        end
        if(_zz_305) begin
          ways_0_metas_45_mru <= 1'b0;
        end
        if(_zz_306) begin
          ways_0_metas_46_mru <= 1'b0;
        end
        if(_zz_307) begin
          ways_0_metas_47_mru <= 1'b0;
        end
        if(_zz_308) begin
          ways_0_metas_48_mru <= 1'b0;
        end
        if(_zz_309) begin
          ways_0_metas_49_mru <= 1'b0;
        end
        if(_zz_310) begin
          ways_0_metas_50_mru <= 1'b0;
        end
        if(_zz_311) begin
          ways_0_metas_51_mru <= 1'b0;
        end
        if(_zz_312) begin
          ways_0_metas_52_mru <= 1'b0;
        end
        if(_zz_313) begin
          ways_0_metas_53_mru <= 1'b0;
        end
        if(_zz_314) begin
          ways_0_metas_54_mru <= 1'b0;
        end
        if(_zz_315) begin
          ways_0_metas_55_mru <= 1'b0;
        end
        if(_zz_316) begin
          ways_0_metas_56_mru <= 1'b0;
        end
        if(_zz_317) begin
          ways_0_metas_57_mru <= 1'b0;
        end
        if(_zz_318) begin
          ways_0_metas_58_mru <= 1'b0;
        end
        if(_zz_319) begin
          ways_0_metas_59_mru <= 1'b0;
        end
        if(_zz_320) begin
          ways_0_metas_60_mru <= 1'b0;
        end
        if(_zz_321) begin
          ways_0_metas_61_mru <= 1'b0;
        end
        if(_zz_322) begin
          ways_0_metas_62_mru <= 1'b0;
        end
        if(_zz_323) begin
          ways_0_metas_63_mru <= 1'b0;
        end
        if(_zz_324) begin
          ways_0_metas_64_mru <= 1'b0;
        end
        if(_zz_325) begin
          ways_0_metas_65_mru <= 1'b0;
        end
        if(_zz_326) begin
          ways_0_metas_66_mru <= 1'b0;
        end
        if(_zz_327) begin
          ways_0_metas_67_mru <= 1'b0;
        end
        if(_zz_328) begin
          ways_0_metas_68_mru <= 1'b0;
        end
        if(_zz_329) begin
          ways_0_metas_69_mru <= 1'b0;
        end
        if(_zz_330) begin
          ways_0_metas_70_mru <= 1'b0;
        end
        if(_zz_331) begin
          ways_0_metas_71_mru <= 1'b0;
        end
        if(_zz_332) begin
          ways_0_metas_72_mru <= 1'b0;
        end
        if(_zz_333) begin
          ways_0_metas_73_mru <= 1'b0;
        end
        if(_zz_334) begin
          ways_0_metas_74_mru <= 1'b0;
        end
        if(_zz_335) begin
          ways_0_metas_75_mru <= 1'b0;
        end
        if(_zz_336) begin
          ways_0_metas_76_mru <= 1'b0;
        end
        if(_zz_337) begin
          ways_0_metas_77_mru <= 1'b0;
        end
        if(_zz_338) begin
          ways_0_metas_78_mru <= 1'b0;
        end
        if(_zz_339) begin
          ways_0_metas_79_mru <= 1'b0;
        end
        if(_zz_340) begin
          ways_0_metas_80_mru <= 1'b0;
        end
        if(_zz_341) begin
          ways_0_metas_81_mru <= 1'b0;
        end
        if(_zz_342) begin
          ways_0_metas_82_mru <= 1'b0;
        end
        if(_zz_343) begin
          ways_0_metas_83_mru <= 1'b0;
        end
        if(_zz_344) begin
          ways_0_metas_84_mru <= 1'b0;
        end
        if(_zz_345) begin
          ways_0_metas_85_mru <= 1'b0;
        end
        if(_zz_346) begin
          ways_0_metas_86_mru <= 1'b0;
        end
        if(_zz_347) begin
          ways_0_metas_87_mru <= 1'b0;
        end
        if(_zz_348) begin
          ways_0_metas_88_mru <= 1'b0;
        end
        if(_zz_349) begin
          ways_0_metas_89_mru <= 1'b0;
        end
        if(_zz_350) begin
          ways_0_metas_90_mru <= 1'b0;
        end
        if(_zz_351) begin
          ways_0_metas_91_mru <= 1'b0;
        end
        if(_zz_352) begin
          ways_0_metas_92_mru <= 1'b0;
        end
        if(_zz_353) begin
          ways_0_metas_93_mru <= 1'b0;
        end
        if(_zz_354) begin
          ways_0_metas_94_mru <= 1'b0;
        end
        if(_zz_355) begin
          ways_0_metas_95_mru <= 1'b0;
        end
        if(_zz_356) begin
          ways_0_metas_96_mru <= 1'b0;
        end
        if(_zz_357) begin
          ways_0_metas_97_mru <= 1'b0;
        end
        if(_zz_358) begin
          ways_0_metas_98_mru <= 1'b0;
        end
        if(_zz_359) begin
          ways_0_metas_99_mru <= 1'b0;
        end
        if(_zz_360) begin
          ways_0_metas_100_mru <= 1'b0;
        end
        if(_zz_361) begin
          ways_0_metas_101_mru <= 1'b0;
        end
        if(_zz_362) begin
          ways_0_metas_102_mru <= 1'b0;
        end
        if(_zz_363) begin
          ways_0_metas_103_mru <= 1'b0;
        end
        if(_zz_364) begin
          ways_0_metas_104_mru <= 1'b0;
        end
        if(_zz_365) begin
          ways_0_metas_105_mru <= 1'b0;
        end
        if(_zz_366) begin
          ways_0_metas_106_mru <= 1'b0;
        end
        if(_zz_367) begin
          ways_0_metas_107_mru <= 1'b0;
        end
        if(_zz_368) begin
          ways_0_metas_108_mru <= 1'b0;
        end
        if(_zz_369) begin
          ways_0_metas_109_mru <= 1'b0;
        end
        if(_zz_370) begin
          ways_0_metas_110_mru <= 1'b0;
        end
        if(_zz_371) begin
          ways_0_metas_111_mru <= 1'b0;
        end
        if(_zz_372) begin
          ways_0_metas_112_mru <= 1'b0;
        end
        if(_zz_373) begin
          ways_0_metas_113_mru <= 1'b0;
        end
        if(_zz_374) begin
          ways_0_metas_114_mru <= 1'b0;
        end
        if(_zz_375) begin
          ways_0_metas_115_mru <= 1'b0;
        end
        if(_zz_376) begin
          ways_0_metas_116_mru <= 1'b0;
        end
        if(_zz_377) begin
          ways_0_metas_117_mru <= 1'b0;
        end
        if(_zz_378) begin
          ways_0_metas_118_mru <= 1'b0;
        end
        if(_zz_379) begin
          ways_0_metas_119_mru <= 1'b0;
        end
        if(_zz_380) begin
          ways_0_metas_120_mru <= 1'b0;
        end
        if(_zz_381) begin
          ways_0_metas_121_mru <= 1'b0;
        end
        if(_zz_382) begin
          ways_0_metas_122_mru <= 1'b0;
        end
        if(_zz_383) begin
          ways_0_metas_123_mru <= 1'b0;
        end
        if(_zz_384) begin
          ways_0_metas_124_mru <= 1'b0;
        end
        if(_zz_385) begin
          ways_0_metas_125_mru <= 1'b0;
        end
        if(_zz_386) begin
          ways_0_metas_126_mru <= 1'b0;
        end
        if(_zz_387) begin
          ways_0_metas_127_mru <= 1'b0;
        end
        if(_zz_260) begin
          ways_0_metas_0_vld <= 1'b0;
        end
        if(_zz_261) begin
          ways_0_metas_1_vld <= 1'b0;
        end
        if(_zz_262) begin
          ways_0_metas_2_vld <= 1'b0;
        end
        if(_zz_263) begin
          ways_0_metas_3_vld <= 1'b0;
        end
        if(_zz_264) begin
          ways_0_metas_4_vld <= 1'b0;
        end
        if(_zz_265) begin
          ways_0_metas_5_vld <= 1'b0;
        end
        if(_zz_266) begin
          ways_0_metas_6_vld <= 1'b0;
        end
        if(_zz_267) begin
          ways_0_metas_7_vld <= 1'b0;
        end
        if(_zz_268) begin
          ways_0_metas_8_vld <= 1'b0;
        end
        if(_zz_269) begin
          ways_0_metas_9_vld <= 1'b0;
        end
        if(_zz_270) begin
          ways_0_metas_10_vld <= 1'b0;
        end
        if(_zz_271) begin
          ways_0_metas_11_vld <= 1'b0;
        end
        if(_zz_272) begin
          ways_0_metas_12_vld <= 1'b0;
        end
        if(_zz_273) begin
          ways_0_metas_13_vld <= 1'b0;
        end
        if(_zz_274) begin
          ways_0_metas_14_vld <= 1'b0;
        end
        if(_zz_275) begin
          ways_0_metas_15_vld <= 1'b0;
        end
        if(_zz_276) begin
          ways_0_metas_16_vld <= 1'b0;
        end
        if(_zz_277) begin
          ways_0_metas_17_vld <= 1'b0;
        end
        if(_zz_278) begin
          ways_0_metas_18_vld <= 1'b0;
        end
        if(_zz_279) begin
          ways_0_metas_19_vld <= 1'b0;
        end
        if(_zz_280) begin
          ways_0_metas_20_vld <= 1'b0;
        end
        if(_zz_281) begin
          ways_0_metas_21_vld <= 1'b0;
        end
        if(_zz_282) begin
          ways_0_metas_22_vld <= 1'b0;
        end
        if(_zz_283) begin
          ways_0_metas_23_vld <= 1'b0;
        end
        if(_zz_284) begin
          ways_0_metas_24_vld <= 1'b0;
        end
        if(_zz_285) begin
          ways_0_metas_25_vld <= 1'b0;
        end
        if(_zz_286) begin
          ways_0_metas_26_vld <= 1'b0;
        end
        if(_zz_287) begin
          ways_0_metas_27_vld <= 1'b0;
        end
        if(_zz_288) begin
          ways_0_metas_28_vld <= 1'b0;
        end
        if(_zz_289) begin
          ways_0_metas_29_vld <= 1'b0;
        end
        if(_zz_290) begin
          ways_0_metas_30_vld <= 1'b0;
        end
        if(_zz_291) begin
          ways_0_metas_31_vld <= 1'b0;
        end
        if(_zz_292) begin
          ways_0_metas_32_vld <= 1'b0;
        end
        if(_zz_293) begin
          ways_0_metas_33_vld <= 1'b0;
        end
        if(_zz_294) begin
          ways_0_metas_34_vld <= 1'b0;
        end
        if(_zz_295) begin
          ways_0_metas_35_vld <= 1'b0;
        end
        if(_zz_296) begin
          ways_0_metas_36_vld <= 1'b0;
        end
        if(_zz_297) begin
          ways_0_metas_37_vld <= 1'b0;
        end
        if(_zz_298) begin
          ways_0_metas_38_vld <= 1'b0;
        end
        if(_zz_299) begin
          ways_0_metas_39_vld <= 1'b0;
        end
        if(_zz_300) begin
          ways_0_metas_40_vld <= 1'b0;
        end
        if(_zz_301) begin
          ways_0_metas_41_vld <= 1'b0;
        end
        if(_zz_302) begin
          ways_0_metas_42_vld <= 1'b0;
        end
        if(_zz_303) begin
          ways_0_metas_43_vld <= 1'b0;
        end
        if(_zz_304) begin
          ways_0_metas_44_vld <= 1'b0;
        end
        if(_zz_305) begin
          ways_0_metas_45_vld <= 1'b0;
        end
        if(_zz_306) begin
          ways_0_metas_46_vld <= 1'b0;
        end
        if(_zz_307) begin
          ways_0_metas_47_vld <= 1'b0;
        end
        if(_zz_308) begin
          ways_0_metas_48_vld <= 1'b0;
        end
        if(_zz_309) begin
          ways_0_metas_49_vld <= 1'b0;
        end
        if(_zz_310) begin
          ways_0_metas_50_vld <= 1'b0;
        end
        if(_zz_311) begin
          ways_0_metas_51_vld <= 1'b0;
        end
        if(_zz_312) begin
          ways_0_metas_52_vld <= 1'b0;
        end
        if(_zz_313) begin
          ways_0_metas_53_vld <= 1'b0;
        end
        if(_zz_314) begin
          ways_0_metas_54_vld <= 1'b0;
        end
        if(_zz_315) begin
          ways_0_metas_55_vld <= 1'b0;
        end
        if(_zz_316) begin
          ways_0_metas_56_vld <= 1'b0;
        end
        if(_zz_317) begin
          ways_0_metas_57_vld <= 1'b0;
        end
        if(_zz_318) begin
          ways_0_metas_58_vld <= 1'b0;
        end
        if(_zz_319) begin
          ways_0_metas_59_vld <= 1'b0;
        end
        if(_zz_320) begin
          ways_0_metas_60_vld <= 1'b0;
        end
        if(_zz_321) begin
          ways_0_metas_61_vld <= 1'b0;
        end
        if(_zz_322) begin
          ways_0_metas_62_vld <= 1'b0;
        end
        if(_zz_323) begin
          ways_0_metas_63_vld <= 1'b0;
        end
        if(_zz_324) begin
          ways_0_metas_64_vld <= 1'b0;
        end
        if(_zz_325) begin
          ways_0_metas_65_vld <= 1'b0;
        end
        if(_zz_326) begin
          ways_0_metas_66_vld <= 1'b0;
        end
        if(_zz_327) begin
          ways_0_metas_67_vld <= 1'b0;
        end
        if(_zz_328) begin
          ways_0_metas_68_vld <= 1'b0;
        end
        if(_zz_329) begin
          ways_0_metas_69_vld <= 1'b0;
        end
        if(_zz_330) begin
          ways_0_metas_70_vld <= 1'b0;
        end
        if(_zz_331) begin
          ways_0_metas_71_vld <= 1'b0;
        end
        if(_zz_332) begin
          ways_0_metas_72_vld <= 1'b0;
        end
        if(_zz_333) begin
          ways_0_metas_73_vld <= 1'b0;
        end
        if(_zz_334) begin
          ways_0_metas_74_vld <= 1'b0;
        end
        if(_zz_335) begin
          ways_0_metas_75_vld <= 1'b0;
        end
        if(_zz_336) begin
          ways_0_metas_76_vld <= 1'b0;
        end
        if(_zz_337) begin
          ways_0_metas_77_vld <= 1'b0;
        end
        if(_zz_338) begin
          ways_0_metas_78_vld <= 1'b0;
        end
        if(_zz_339) begin
          ways_0_metas_79_vld <= 1'b0;
        end
        if(_zz_340) begin
          ways_0_metas_80_vld <= 1'b0;
        end
        if(_zz_341) begin
          ways_0_metas_81_vld <= 1'b0;
        end
        if(_zz_342) begin
          ways_0_metas_82_vld <= 1'b0;
        end
        if(_zz_343) begin
          ways_0_metas_83_vld <= 1'b0;
        end
        if(_zz_344) begin
          ways_0_metas_84_vld <= 1'b0;
        end
        if(_zz_345) begin
          ways_0_metas_85_vld <= 1'b0;
        end
        if(_zz_346) begin
          ways_0_metas_86_vld <= 1'b0;
        end
        if(_zz_347) begin
          ways_0_metas_87_vld <= 1'b0;
        end
        if(_zz_348) begin
          ways_0_metas_88_vld <= 1'b0;
        end
        if(_zz_349) begin
          ways_0_metas_89_vld <= 1'b0;
        end
        if(_zz_350) begin
          ways_0_metas_90_vld <= 1'b0;
        end
        if(_zz_351) begin
          ways_0_metas_91_vld <= 1'b0;
        end
        if(_zz_352) begin
          ways_0_metas_92_vld <= 1'b0;
        end
        if(_zz_353) begin
          ways_0_metas_93_vld <= 1'b0;
        end
        if(_zz_354) begin
          ways_0_metas_94_vld <= 1'b0;
        end
        if(_zz_355) begin
          ways_0_metas_95_vld <= 1'b0;
        end
        if(_zz_356) begin
          ways_0_metas_96_vld <= 1'b0;
        end
        if(_zz_357) begin
          ways_0_metas_97_vld <= 1'b0;
        end
        if(_zz_358) begin
          ways_0_metas_98_vld <= 1'b0;
        end
        if(_zz_359) begin
          ways_0_metas_99_vld <= 1'b0;
        end
        if(_zz_360) begin
          ways_0_metas_100_vld <= 1'b0;
        end
        if(_zz_361) begin
          ways_0_metas_101_vld <= 1'b0;
        end
        if(_zz_362) begin
          ways_0_metas_102_vld <= 1'b0;
        end
        if(_zz_363) begin
          ways_0_metas_103_vld <= 1'b0;
        end
        if(_zz_364) begin
          ways_0_metas_104_vld <= 1'b0;
        end
        if(_zz_365) begin
          ways_0_metas_105_vld <= 1'b0;
        end
        if(_zz_366) begin
          ways_0_metas_106_vld <= 1'b0;
        end
        if(_zz_367) begin
          ways_0_metas_107_vld <= 1'b0;
        end
        if(_zz_368) begin
          ways_0_metas_108_vld <= 1'b0;
        end
        if(_zz_369) begin
          ways_0_metas_109_vld <= 1'b0;
        end
        if(_zz_370) begin
          ways_0_metas_110_vld <= 1'b0;
        end
        if(_zz_371) begin
          ways_0_metas_111_vld <= 1'b0;
        end
        if(_zz_372) begin
          ways_0_metas_112_vld <= 1'b0;
        end
        if(_zz_373) begin
          ways_0_metas_113_vld <= 1'b0;
        end
        if(_zz_374) begin
          ways_0_metas_114_vld <= 1'b0;
        end
        if(_zz_375) begin
          ways_0_metas_115_vld <= 1'b0;
        end
        if(_zz_376) begin
          ways_0_metas_116_vld <= 1'b0;
        end
        if(_zz_377) begin
          ways_0_metas_117_vld <= 1'b0;
        end
        if(_zz_378) begin
          ways_0_metas_118_vld <= 1'b0;
        end
        if(_zz_379) begin
          ways_0_metas_119_vld <= 1'b0;
        end
        if(_zz_380) begin
          ways_0_metas_120_vld <= 1'b0;
        end
        if(_zz_381) begin
          ways_0_metas_121_vld <= 1'b0;
        end
        if(_zz_382) begin
          ways_0_metas_122_vld <= 1'b0;
        end
        if(_zz_383) begin
          ways_0_metas_123_vld <= 1'b0;
        end
        if(_zz_384) begin
          ways_0_metas_124_vld <= 1'b0;
        end
        if(_zz_385) begin
          ways_0_metas_125_vld <= 1'b0;
        end
        if(_zz_386) begin
          ways_0_metas_126_vld <= 1'b0;
        end
        if(_zz_387) begin
          ways_0_metas_127_vld <= 1'b0;
        end
      end else begin
        if(when_ICache_l210) begin
          if(cache_hit_0) begin
            if(_zz_2) begin
              ways_0_metas_0_mru <= 1'b1;
            end
            if(_zz_3) begin
              ways_0_metas_1_mru <= 1'b1;
            end
            if(_zz_4) begin
              ways_0_metas_2_mru <= 1'b1;
            end
            if(_zz_5) begin
              ways_0_metas_3_mru <= 1'b1;
            end
            if(_zz_6) begin
              ways_0_metas_4_mru <= 1'b1;
            end
            if(_zz_7) begin
              ways_0_metas_5_mru <= 1'b1;
            end
            if(_zz_8) begin
              ways_0_metas_6_mru <= 1'b1;
            end
            if(_zz_9) begin
              ways_0_metas_7_mru <= 1'b1;
            end
            if(_zz_10) begin
              ways_0_metas_8_mru <= 1'b1;
            end
            if(_zz_11) begin
              ways_0_metas_9_mru <= 1'b1;
            end
            if(_zz_12) begin
              ways_0_metas_10_mru <= 1'b1;
            end
            if(_zz_13) begin
              ways_0_metas_11_mru <= 1'b1;
            end
            if(_zz_14) begin
              ways_0_metas_12_mru <= 1'b1;
            end
            if(_zz_15) begin
              ways_0_metas_13_mru <= 1'b1;
            end
            if(_zz_16) begin
              ways_0_metas_14_mru <= 1'b1;
            end
            if(_zz_17) begin
              ways_0_metas_15_mru <= 1'b1;
            end
            if(_zz_18) begin
              ways_0_metas_16_mru <= 1'b1;
            end
            if(_zz_19) begin
              ways_0_metas_17_mru <= 1'b1;
            end
            if(_zz_20) begin
              ways_0_metas_18_mru <= 1'b1;
            end
            if(_zz_21) begin
              ways_0_metas_19_mru <= 1'b1;
            end
            if(_zz_22) begin
              ways_0_metas_20_mru <= 1'b1;
            end
            if(_zz_23) begin
              ways_0_metas_21_mru <= 1'b1;
            end
            if(_zz_24) begin
              ways_0_metas_22_mru <= 1'b1;
            end
            if(_zz_25) begin
              ways_0_metas_23_mru <= 1'b1;
            end
            if(_zz_26) begin
              ways_0_metas_24_mru <= 1'b1;
            end
            if(_zz_27) begin
              ways_0_metas_25_mru <= 1'b1;
            end
            if(_zz_28) begin
              ways_0_metas_26_mru <= 1'b1;
            end
            if(_zz_29) begin
              ways_0_metas_27_mru <= 1'b1;
            end
            if(_zz_30) begin
              ways_0_metas_28_mru <= 1'b1;
            end
            if(_zz_31) begin
              ways_0_metas_29_mru <= 1'b1;
            end
            if(_zz_32) begin
              ways_0_metas_30_mru <= 1'b1;
            end
            if(_zz_33) begin
              ways_0_metas_31_mru <= 1'b1;
            end
            if(_zz_34) begin
              ways_0_metas_32_mru <= 1'b1;
            end
            if(_zz_35) begin
              ways_0_metas_33_mru <= 1'b1;
            end
            if(_zz_36) begin
              ways_0_metas_34_mru <= 1'b1;
            end
            if(_zz_37) begin
              ways_0_metas_35_mru <= 1'b1;
            end
            if(_zz_38) begin
              ways_0_metas_36_mru <= 1'b1;
            end
            if(_zz_39) begin
              ways_0_metas_37_mru <= 1'b1;
            end
            if(_zz_40) begin
              ways_0_metas_38_mru <= 1'b1;
            end
            if(_zz_41) begin
              ways_0_metas_39_mru <= 1'b1;
            end
            if(_zz_42) begin
              ways_0_metas_40_mru <= 1'b1;
            end
            if(_zz_43) begin
              ways_0_metas_41_mru <= 1'b1;
            end
            if(_zz_44) begin
              ways_0_metas_42_mru <= 1'b1;
            end
            if(_zz_45) begin
              ways_0_metas_43_mru <= 1'b1;
            end
            if(_zz_46) begin
              ways_0_metas_44_mru <= 1'b1;
            end
            if(_zz_47) begin
              ways_0_metas_45_mru <= 1'b1;
            end
            if(_zz_48) begin
              ways_0_metas_46_mru <= 1'b1;
            end
            if(_zz_49) begin
              ways_0_metas_47_mru <= 1'b1;
            end
            if(_zz_50) begin
              ways_0_metas_48_mru <= 1'b1;
            end
            if(_zz_51) begin
              ways_0_metas_49_mru <= 1'b1;
            end
            if(_zz_52) begin
              ways_0_metas_50_mru <= 1'b1;
            end
            if(_zz_53) begin
              ways_0_metas_51_mru <= 1'b1;
            end
            if(_zz_54) begin
              ways_0_metas_52_mru <= 1'b1;
            end
            if(_zz_55) begin
              ways_0_metas_53_mru <= 1'b1;
            end
            if(_zz_56) begin
              ways_0_metas_54_mru <= 1'b1;
            end
            if(_zz_57) begin
              ways_0_metas_55_mru <= 1'b1;
            end
            if(_zz_58) begin
              ways_0_metas_56_mru <= 1'b1;
            end
            if(_zz_59) begin
              ways_0_metas_57_mru <= 1'b1;
            end
            if(_zz_60) begin
              ways_0_metas_58_mru <= 1'b1;
            end
            if(_zz_61) begin
              ways_0_metas_59_mru <= 1'b1;
            end
            if(_zz_62) begin
              ways_0_metas_60_mru <= 1'b1;
            end
            if(_zz_63) begin
              ways_0_metas_61_mru <= 1'b1;
            end
            if(_zz_64) begin
              ways_0_metas_62_mru <= 1'b1;
            end
            if(_zz_65) begin
              ways_0_metas_63_mru <= 1'b1;
            end
            if(_zz_66) begin
              ways_0_metas_64_mru <= 1'b1;
            end
            if(_zz_67) begin
              ways_0_metas_65_mru <= 1'b1;
            end
            if(_zz_68) begin
              ways_0_metas_66_mru <= 1'b1;
            end
            if(_zz_69) begin
              ways_0_metas_67_mru <= 1'b1;
            end
            if(_zz_70) begin
              ways_0_metas_68_mru <= 1'b1;
            end
            if(_zz_71) begin
              ways_0_metas_69_mru <= 1'b1;
            end
            if(_zz_72) begin
              ways_0_metas_70_mru <= 1'b1;
            end
            if(_zz_73) begin
              ways_0_metas_71_mru <= 1'b1;
            end
            if(_zz_74) begin
              ways_0_metas_72_mru <= 1'b1;
            end
            if(_zz_75) begin
              ways_0_metas_73_mru <= 1'b1;
            end
            if(_zz_76) begin
              ways_0_metas_74_mru <= 1'b1;
            end
            if(_zz_77) begin
              ways_0_metas_75_mru <= 1'b1;
            end
            if(_zz_78) begin
              ways_0_metas_76_mru <= 1'b1;
            end
            if(_zz_79) begin
              ways_0_metas_77_mru <= 1'b1;
            end
            if(_zz_80) begin
              ways_0_metas_78_mru <= 1'b1;
            end
            if(_zz_81) begin
              ways_0_metas_79_mru <= 1'b1;
            end
            if(_zz_82) begin
              ways_0_metas_80_mru <= 1'b1;
            end
            if(_zz_83) begin
              ways_0_metas_81_mru <= 1'b1;
            end
            if(_zz_84) begin
              ways_0_metas_82_mru <= 1'b1;
            end
            if(_zz_85) begin
              ways_0_metas_83_mru <= 1'b1;
            end
            if(_zz_86) begin
              ways_0_metas_84_mru <= 1'b1;
            end
            if(_zz_87) begin
              ways_0_metas_85_mru <= 1'b1;
            end
            if(_zz_88) begin
              ways_0_metas_86_mru <= 1'b1;
            end
            if(_zz_89) begin
              ways_0_metas_87_mru <= 1'b1;
            end
            if(_zz_90) begin
              ways_0_metas_88_mru <= 1'b1;
            end
            if(_zz_91) begin
              ways_0_metas_89_mru <= 1'b1;
            end
            if(_zz_92) begin
              ways_0_metas_90_mru <= 1'b1;
            end
            if(_zz_93) begin
              ways_0_metas_91_mru <= 1'b1;
            end
            if(_zz_94) begin
              ways_0_metas_92_mru <= 1'b1;
            end
            if(_zz_95) begin
              ways_0_metas_93_mru <= 1'b1;
            end
            if(_zz_96) begin
              ways_0_metas_94_mru <= 1'b1;
            end
            if(_zz_97) begin
              ways_0_metas_95_mru <= 1'b1;
            end
            if(_zz_98) begin
              ways_0_metas_96_mru <= 1'b1;
            end
            if(_zz_99) begin
              ways_0_metas_97_mru <= 1'b1;
            end
            if(_zz_100) begin
              ways_0_metas_98_mru <= 1'b1;
            end
            if(_zz_101) begin
              ways_0_metas_99_mru <= 1'b1;
            end
            if(_zz_102) begin
              ways_0_metas_100_mru <= 1'b1;
            end
            if(_zz_103) begin
              ways_0_metas_101_mru <= 1'b1;
            end
            if(_zz_104) begin
              ways_0_metas_102_mru <= 1'b1;
            end
            if(_zz_105) begin
              ways_0_metas_103_mru <= 1'b1;
            end
            if(_zz_106) begin
              ways_0_metas_104_mru <= 1'b1;
            end
            if(_zz_107) begin
              ways_0_metas_105_mru <= 1'b1;
            end
            if(_zz_108) begin
              ways_0_metas_106_mru <= 1'b1;
            end
            if(_zz_109) begin
              ways_0_metas_107_mru <= 1'b1;
            end
            if(_zz_110) begin
              ways_0_metas_108_mru <= 1'b1;
            end
            if(_zz_111) begin
              ways_0_metas_109_mru <= 1'b1;
            end
            if(_zz_112) begin
              ways_0_metas_110_mru <= 1'b1;
            end
            if(_zz_113) begin
              ways_0_metas_111_mru <= 1'b1;
            end
            if(_zz_114) begin
              ways_0_metas_112_mru <= 1'b1;
            end
            if(_zz_115) begin
              ways_0_metas_113_mru <= 1'b1;
            end
            if(_zz_116) begin
              ways_0_metas_114_mru <= 1'b1;
            end
            if(_zz_117) begin
              ways_0_metas_115_mru <= 1'b1;
            end
            if(_zz_118) begin
              ways_0_metas_116_mru <= 1'b1;
            end
            if(_zz_119) begin
              ways_0_metas_117_mru <= 1'b1;
            end
            if(_zz_120) begin
              ways_0_metas_118_mru <= 1'b1;
            end
            if(_zz_121) begin
              ways_0_metas_119_mru <= 1'b1;
            end
            if(_zz_122) begin
              ways_0_metas_120_mru <= 1'b1;
            end
            if(_zz_123) begin
              ways_0_metas_121_mru <= 1'b1;
            end
            if(_zz_124) begin
              ways_0_metas_122_mru <= 1'b1;
            end
            if(_zz_125) begin
              ways_0_metas_123_mru <= 1'b1;
            end
            if(_zz_126) begin
              ways_0_metas_124_mru <= 1'b1;
            end
            if(_zz_127) begin
              ways_0_metas_125_mru <= 1'b1;
            end
            if(_zz_128) begin
              ways_0_metas_126_mru <= 1'b1;
            end
            if(_zz_129) begin
              ways_0_metas_127_mru <= 1'b1;
            end
          end else begin
            if(_zz_2) begin
              ways_0_metas_0_mru <= 1'b0;
            end
            if(_zz_3) begin
              ways_0_metas_1_mru <= 1'b0;
            end
            if(_zz_4) begin
              ways_0_metas_2_mru <= 1'b0;
            end
            if(_zz_5) begin
              ways_0_metas_3_mru <= 1'b0;
            end
            if(_zz_6) begin
              ways_0_metas_4_mru <= 1'b0;
            end
            if(_zz_7) begin
              ways_0_metas_5_mru <= 1'b0;
            end
            if(_zz_8) begin
              ways_0_metas_6_mru <= 1'b0;
            end
            if(_zz_9) begin
              ways_0_metas_7_mru <= 1'b0;
            end
            if(_zz_10) begin
              ways_0_metas_8_mru <= 1'b0;
            end
            if(_zz_11) begin
              ways_0_metas_9_mru <= 1'b0;
            end
            if(_zz_12) begin
              ways_0_metas_10_mru <= 1'b0;
            end
            if(_zz_13) begin
              ways_0_metas_11_mru <= 1'b0;
            end
            if(_zz_14) begin
              ways_0_metas_12_mru <= 1'b0;
            end
            if(_zz_15) begin
              ways_0_metas_13_mru <= 1'b0;
            end
            if(_zz_16) begin
              ways_0_metas_14_mru <= 1'b0;
            end
            if(_zz_17) begin
              ways_0_metas_15_mru <= 1'b0;
            end
            if(_zz_18) begin
              ways_0_metas_16_mru <= 1'b0;
            end
            if(_zz_19) begin
              ways_0_metas_17_mru <= 1'b0;
            end
            if(_zz_20) begin
              ways_0_metas_18_mru <= 1'b0;
            end
            if(_zz_21) begin
              ways_0_metas_19_mru <= 1'b0;
            end
            if(_zz_22) begin
              ways_0_metas_20_mru <= 1'b0;
            end
            if(_zz_23) begin
              ways_0_metas_21_mru <= 1'b0;
            end
            if(_zz_24) begin
              ways_0_metas_22_mru <= 1'b0;
            end
            if(_zz_25) begin
              ways_0_metas_23_mru <= 1'b0;
            end
            if(_zz_26) begin
              ways_0_metas_24_mru <= 1'b0;
            end
            if(_zz_27) begin
              ways_0_metas_25_mru <= 1'b0;
            end
            if(_zz_28) begin
              ways_0_metas_26_mru <= 1'b0;
            end
            if(_zz_29) begin
              ways_0_metas_27_mru <= 1'b0;
            end
            if(_zz_30) begin
              ways_0_metas_28_mru <= 1'b0;
            end
            if(_zz_31) begin
              ways_0_metas_29_mru <= 1'b0;
            end
            if(_zz_32) begin
              ways_0_metas_30_mru <= 1'b0;
            end
            if(_zz_33) begin
              ways_0_metas_31_mru <= 1'b0;
            end
            if(_zz_34) begin
              ways_0_metas_32_mru <= 1'b0;
            end
            if(_zz_35) begin
              ways_0_metas_33_mru <= 1'b0;
            end
            if(_zz_36) begin
              ways_0_metas_34_mru <= 1'b0;
            end
            if(_zz_37) begin
              ways_0_metas_35_mru <= 1'b0;
            end
            if(_zz_38) begin
              ways_0_metas_36_mru <= 1'b0;
            end
            if(_zz_39) begin
              ways_0_metas_37_mru <= 1'b0;
            end
            if(_zz_40) begin
              ways_0_metas_38_mru <= 1'b0;
            end
            if(_zz_41) begin
              ways_0_metas_39_mru <= 1'b0;
            end
            if(_zz_42) begin
              ways_0_metas_40_mru <= 1'b0;
            end
            if(_zz_43) begin
              ways_0_metas_41_mru <= 1'b0;
            end
            if(_zz_44) begin
              ways_0_metas_42_mru <= 1'b0;
            end
            if(_zz_45) begin
              ways_0_metas_43_mru <= 1'b0;
            end
            if(_zz_46) begin
              ways_0_metas_44_mru <= 1'b0;
            end
            if(_zz_47) begin
              ways_0_metas_45_mru <= 1'b0;
            end
            if(_zz_48) begin
              ways_0_metas_46_mru <= 1'b0;
            end
            if(_zz_49) begin
              ways_0_metas_47_mru <= 1'b0;
            end
            if(_zz_50) begin
              ways_0_metas_48_mru <= 1'b0;
            end
            if(_zz_51) begin
              ways_0_metas_49_mru <= 1'b0;
            end
            if(_zz_52) begin
              ways_0_metas_50_mru <= 1'b0;
            end
            if(_zz_53) begin
              ways_0_metas_51_mru <= 1'b0;
            end
            if(_zz_54) begin
              ways_0_metas_52_mru <= 1'b0;
            end
            if(_zz_55) begin
              ways_0_metas_53_mru <= 1'b0;
            end
            if(_zz_56) begin
              ways_0_metas_54_mru <= 1'b0;
            end
            if(_zz_57) begin
              ways_0_metas_55_mru <= 1'b0;
            end
            if(_zz_58) begin
              ways_0_metas_56_mru <= 1'b0;
            end
            if(_zz_59) begin
              ways_0_metas_57_mru <= 1'b0;
            end
            if(_zz_60) begin
              ways_0_metas_58_mru <= 1'b0;
            end
            if(_zz_61) begin
              ways_0_metas_59_mru <= 1'b0;
            end
            if(_zz_62) begin
              ways_0_metas_60_mru <= 1'b0;
            end
            if(_zz_63) begin
              ways_0_metas_61_mru <= 1'b0;
            end
            if(_zz_64) begin
              ways_0_metas_62_mru <= 1'b0;
            end
            if(_zz_65) begin
              ways_0_metas_63_mru <= 1'b0;
            end
            if(_zz_66) begin
              ways_0_metas_64_mru <= 1'b0;
            end
            if(_zz_67) begin
              ways_0_metas_65_mru <= 1'b0;
            end
            if(_zz_68) begin
              ways_0_metas_66_mru <= 1'b0;
            end
            if(_zz_69) begin
              ways_0_metas_67_mru <= 1'b0;
            end
            if(_zz_70) begin
              ways_0_metas_68_mru <= 1'b0;
            end
            if(_zz_71) begin
              ways_0_metas_69_mru <= 1'b0;
            end
            if(_zz_72) begin
              ways_0_metas_70_mru <= 1'b0;
            end
            if(_zz_73) begin
              ways_0_metas_71_mru <= 1'b0;
            end
            if(_zz_74) begin
              ways_0_metas_72_mru <= 1'b0;
            end
            if(_zz_75) begin
              ways_0_metas_73_mru <= 1'b0;
            end
            if(_zz_76) begin
              ways_0_metas_74_mru <= 1'b0;
            end
            if(_zz_77) begin
              ways_0_metas_75_mru <= 1'b0;
            end
            if(_zz_78) begin
              ways_0_metas_76_mru <= 1'b0;
            end
            if(_zz_79) begin
              ways_0_metas_77_mru <= 1'b0;
            end
            if(_zz_80) begin
              ways_0_metas_78_mru <= 1'b0;
            end
            if(_zz_81) begin
              ways_0_metas_79_mru <= 1'b0;
            end
            if(_zz_82) begin
              ways_0_metas_80_mru <= 1'b0;
            end
            if(_zz_83) begin
              ways_0_metas_81_mru <= 1'b0;
            end
            if(_zz_84) begin
              ways_0_metas_82_mru <= 1'b0;
            end
            if(_zz_85) begin
              ways_0_metas_83_mru <= 1'b0;
            end
            if(_zz_86) begin
              ways_0_metas_84_mru <= 1'b0;
            end
            if(_zz_87) begin
              ways_0_metas_85_mru <= 1'b0;
            end
            if(_zz_88) begin
              ways_0_metas_86_mru <= 1'b0;
            end
            if(_zz_89) begin
              ways_0_metas_87_mru <= 1'b0;
            end
            if(_zz_90) begin
              ways_0_metas_88_mru <= 1'b0;
            end
            if(_zz_91) begin
              ways_0_metas_89_mru <= 1'b0;
            end
            if(_zz_92) begin
              ways_0_metas_90_mru <= 1'b0;
            end
            if(_zz_93) begin
              ways_0_metas_91_mru <= 1'b0;
            end
            if(_zz_94) begin
              ways_0_metas_92_mru <= 1'b0;
            end
            if(_zz_95) begin
              ways_0_metas_93_mru <= 1'b0;
            end
            if(_zz_96) begin
              ways_0_metas_94_mru <= 1'b0;
            end
            if(_zz_97) begin
              ways_0_metas_95_mru <= 1'b0;
            end
            if(_zz_98) begin
              ways_0_metas_96_mru <= 1'b0;
            end
            if(_zz_99) begin
              ways_0_metas_97_mru <= 1'b0;
            end
            if(_zz_100) begin
              ways_0_metas_98_mru <= 1'b0;
            end
            if(_zz_101) begin
              ways_0_metas_99_mru <= 1'b0;
            end
            if(_zz_102) begin
              ways_0_metas_100_mru <= 1'b0;
            end
            if(_zz_103) begin
              ways_0_metas_101_mru <= 1'b0;
            end
            if(_zz_104) begin
              ways_0_metas_102_mru <= 1'b0;
            end
            if(_zz_105) begin
              ways_0_metas_103_mru <= 1'b0;
            end
            if(_zz_106) begin
              ways_0_metas_104_mru <= 1'b0;
            end
            if(_zz_107) begin
              ways_0_metas_105_mru <= 1'b0;
            end
            if(_zz_108) begin
              ways_0_metas_106_mru <= 1'b0;
            end
            if(_zz_109) begin
              ways_0_metas_107_mru <= 1'b0;
            end
            if(_zz_110) begin
              ways_0_metas_108_mru <= 1'b0;
            end
            if(_zz_111) begin
              ways_0_metas_109_mru <= 1'b0;
            end
            if(_zz_112) begin
              ways_0_metas_110_mru <= 1'b0;
            end
            if(_zz_113) begin
              ways_0_metas_111_mru <= 1'b0;
            end
            if(_zz_114) begin
              ways_0_metas_112_mru <= 1'b0;
            end
            if(_zz_115) begin
              ways_0_metas_113_mru <= 1'b0;
            end
            if(_zz_116) begin
              ways_0_metas_114_mru <= 1'b0;
            end
            if(_zz_117) begin
              ways_0_metas_115_mru <= 1'b0;
            end
            if(_zz_118) begin
              ways_0_metas_116_mru <= 1'b0;
            end
            if(_zz_119) begin
              ways_0_metas_117_mru <= 1'b0;
            end
            if(_zz_120) begin
              ways_0_metas_118_mru <= 1'b0;
            end
            if(_zz_121) begin
              ways_0_metas_119_mru <= 1'b0;
            end
            if(_zz_122) begin
              ways_0_metas_120_mru <= 1'b0;
            end
            if(_zz_123) begin
              ways_0_metas_121_mru <= 1'b0;
            end
            if(_zz_124) begin
              ways_0_metas_122_mru <= 1'b0;
            end
            if(_zz_125) begin
              ways_0_metas_123_mru <= 1'b0;
            end
            if(_zz_126) begin
              ways_0_metas_124_mru <= 1'b0;
            end
            if(_zz_127) begin
              ways_0_metas_125_mru <= 1'b0;
            end
            if(_zz_128) begin
              ways_0_metas_126_mru <= 1'b0;
            end
            if(_zz_129) begin
              ways_0_metas_127_mru <= 1'b0;
            end
          end
        end else begin
          if(when_ICache_l217) begin
            if(_zz_2) begin
              ways_0_metas_0_mru <= 1'b1;
            end
            if(_zz_3) begin
              ways_0_metas_1_mru <= 1'b1;
            end
            if(_zz_4) begin
              ways_0_metas_2_mru <= 1'b1;
            end
            if(_zz_5) begin
              ways_0_metas_3_mru <= 1'b1;
            end
            if(_zz_6) begin
              ways_0_metas_4_mru <= 1'b1;
            end
            if(_zz_7) begin
              ways_0_metas_5_mru <= 1'b1;
            end
            if(_zz_8) begin
              ways_0_metas_6_mru <= 1'b1;
            end
            if(_zz_9) begin
              ways_0_metas_7_mru <= 1'b1;
            end
            if(_zz_10) begin
              ways_0_metas_8_mru <= 1'b1;
            end
            if(_zz_11) begin
              ways_0_metas_9_mru <= 1'b1;
            end
            if(_zz_12) begin
              ways_0_metas_10_mru <= 1'b1;
            end
            if(_zz_13) begin
              ways_0_metas_11_mru <= 1'b1;
            end
            if(_zz_14) begin
              ways_0_metas_12_mru <= 1'b1;
            end
            if(_zz_15) begin
              ways_0_metas_13_mru <= 1'b1;
            end
            if(_zz_16) begin
              ways_0_metas_14_mru <= 1'b1;
            end
            if(_zz_17) begin
              ways_0_metas_15_mru <= 1'b1;
            end
            if(_zz_18) begin
              ways_0_metas_16_mru <= 1'b1;
            end
            if(_zz_19) begin
              ways_0_metas_17_mru <= 1'b1;
            end
            if(_zz_20) begin
              ways_0_metas_18_mru <= 1'b1;
            end
            if(_zz_21) begin
              ways_0_metas_19_mru <= 1'b1;
            end
            if(_zz_22) begin
              ways_0_metas_20_mru <= 1'b1;
            end
            if(_zz_23) begin
              ways_0_metas_21_mru <= 1'b1;
            end
            if(_zz_24) begin
              ways_0_metas_22_mru <= 1'b1;
            end
            if(_zz_25) begin
              ways_0_metas_23_mru <= 1'b1;
            end
            if(_zz_26) begin
              ways_0_metas_24_mru <= 1'b1;
            end
            if(_zz_27) begin
              ways_0_metas_25_mru <= 1'b1;
            end
            if(_zz_28) begin
              ways_0_metas_26_mru <= 1'b1;
            end
            if(_zz_29) begin
              ways_0_metas_27_mru <= 1'b1;
            end
            if(_zz_30) begin
              ways_0_metas_28_mru <= 1'b1;
            end
            if(_zz_31) begin
              ways_0_metas_29_mru <= 1'b1;
            end
            if(_zz_32) begin
              ways_0_metas_30_mru <= 1'b1;
            end
            if(_zz_33) begin
              ways_0_metas_31_mru <= 1'b1;
            end
            if(_zz_34) begin
              ways_0_metas_32_mru <= 1'b1;
            end
            if(_zz_35) begin
              ways_0_metas_33_mru <= 1'b1;
            end
            if(_zz_36) begin
              ways_0_metas_34_mru <= 1'b1;
            end
            if(_zz_37) begin
              ways_0_metas_35_mru <= 1'b1;
            end
            if(_zz_38) begin
              ways_0_metas_36_mru <= 1'b1;
            end
            if(_zz_39) begin
              ways_0_metas_37_mru <= 1'b1;
            end
            if(_zz_40) begin
              ways_0_metas_38_mru <= 1'b1;
            end
            if(_zz_41) begin
              ways_0_metas_39_mru <= 1'b1;
            end
            if(_zz_42) begin
              ways_0_metas_40_mru <= 1'b1;
            end
            if(_zz_43) begin
              ways_0_metas_41_mru <= 1'b1;
            end
            if(_zz_44) begin
              ways_0_metas_42_mru <= 1'b1;
            end
            if(_zz_45) begin
              ways_0_metas_43_mru <= 1'b1;
            end
            if(_zz_46) begin
              ways_0_metas_44_mru <= 1'b1;
            end
            if(_zz_47) begin
              ways_0_metas_45_mru <= 1'b1;
            end
            if(_zz_48) begin
              ways_0_metas_46_mru <= 1'b1;
            end
            if(_zz_49) begin
              ways_0_metas_47_mru <= 1'b1;
            end
            if(_zz_50) begin
              ways_0_metas_48_mru <= 1'b1;
            end
            if(_zz_51) begin
              ways_0_metas_49_mru <= 1'b1;
            end
            if(_zz_52) begin
              ways_0_metas_50_mru <= 1'b1;
            end
            if(_zz_53) begin
              ways_0_metas_51_mru <= 1'b1;
            end
            if(_zz_54) begin
              ways_0_metas_52_mru <= 1'b1;
            end
            if(_zz_55) begin
              ways_0_metas_53_mru <= 1'b1;
            end
            if(_zz_56) begin
              ways_0_metas_54_mru <= 1'b1;
            end
            if(_zz_57) begin
              ways_0_metas_55_mru <= 1'b1;
            end
            if(_zz_58) begin
              ways_0_metas_56_mru <= 1'b1;
            end
            if(_zz_59) begin
              ways_0_metas_57_mru <= 1'b1;
            end
            if(_zz_60) begin
              ways_0_metas_58_mru <= 1'b1;
            end
            if(_zz_61) begin
              ways_0_metas_59_mru <= 1'b1;
            end
            if(_zz_62) begin
              ways_0_metas_60_mru <= 1'b1;
            end
            if(_zz_63) begin
              ways_0_metas_61_mru <= 1'b1;
            end
            if(_zz_64) begin
              ways_0_metas_62_mru <= 1'b1;
            end
            if(_zz_65) begin
              ways_0_metas_63_mru <= 1'b1;
            end
            if(_zz_66) begin
              ways_0_metas_64_mru <= 1'b1;
            end
            if(_zz_67) begin
              ways_0_metas_65_mru <= 1'b1;
            end
            if(_zz_68) begin
              ways_0_metas_66_mru <= 1'b1;
            end
            if(_zz_69) begin
              ways_0_metas_67_mru <= 1'b1;
            end
            if(_zz_70) begin
              ways_0_metas_68_mru <= 1'b1;
            end
            if(_zz_71) begin
              ways_0_metas_69_mru <= 1'b1;
            end
            if(_zz_72) begin
              ways_0_metas_70_mru <= 1'b1;
            end
            if(_zz_73) begin
              ways_0_metas_71_mru <= 1'b1;
            end
            if(_zz_74) begin
              ways_0_metas_72_mru <= 1'b1;
            end
            if(_zz_75) begin
              ways_0_metas_73_mru <= 1'b1;
            end
            if(_zz_76) begin
              ways_0_metas_74_mru <= 1'b1;
            end
            if(_zz_77) begin
              ways_0_metas_75_mru <= 1'b1;
            end
            if(_zz_78) begin
              ways_0_metas_76_mru <= 1'b1;
            end
            if(_zz_79) begin
              ways_0_metas_77_mru <= 1'b1;
            end
            if(_zz_80) begin
              ways_0_metas_78_mru <= 1'b1;
            end
            if(_zz_81) begin
              ways_0_metas_79_mru <= 1'b1;
            end
            if(_zz_82) begin
              ways_0_metas_80_mru <= 1'b1;
            end
            if(_zz_83) begin
              ways_0_metas_81_mru <= 1'b1;
            end
            if(_zz_84) begin
              ways_0_metas_82_mru <= 1'b1;
            end
            if(_zz_85) begin
              ways_0_metas_83_mru <= 1'b1;
            end
            if(_zz_86) begin
              ways_0_metas_84_mru <= 1'b1;
            end
            if(_zz_87) begin
              ways_0_metas_85_mru <= 1'b1;
            end
            if(_zz_88) begin
              ways_0_metas_86_mru <= 1'b1;
            end
            if(_zz_89) begin
              ways_0_metas_87_mru <= 1'b1;
            end
            if(_zz_90) begin
              ways_0_metas_88_mru <= 1'b1;
            end
            if(_zz_91) begin
              ways_0_metas_89_mru <= 1'b1;
            end
            if(_zz_92) begin
              ways_0_metas_90_mru <= 1'b1;
            end
            if(_zz_93) begin
              ways_0_metas_91_mru <= 1'b1;
            end
            if(_zz_94) begin
              ways_0_metas_92_mru <= 1'b1;
            end
            if(_zz_95) begin
              ways_0_metas_93_mru <= 1'b1;
            end
            if(_zz_96) begin
              ways_0_metas_94_mru <= 1'b1;
            end
            if(_zz_97) begin
              ways_0_metas_95_mru <= 1'b1;
            end
            if(_zz_98) begin
              ways_0_metas_96_mru <= 1'b1;
            end
            if(_zz_99) begin
              ways_0_metas_97_mru <= 1'b1;
            end
            if(_zz_100) begin
              ways_0_metas_98_mru <= 1'b1;
            end
            if(_zz_101) begin
              ways_0_metas_99_mru <= 1'b1;
            end
            if(_zz_102) begin
              ways_0_metas_100_mru <= 1'b1;
            end
            if(_zz_103) begin
              ways_0_metas_101_mru <= 1'b1;
            end
            if(_zz_104) begin
              ways_0_metas_102_mru <= 1'b1;
            end
            if(_zz_105) begin
              ways_0_metas_103_mru <= 1'b1;
            end
            if(_zz_106) begin
              ways_0_metas_104_mru <= 1'b1;
            end
            if(_zz_107) begin
              ways_0_metas_105_mru <= 1'b1;
            end
            if(_zz_108) begin
              ways_0_metas_106_mru <= 1'b1;
            end
            if(_zz_109) begin
              ways_0_metas_107_mru <= 1'b1;
            end
            if(_zz_110) begin
              ways_0_metas_108_mru <= 1'b1;
            end
            if(_zz_111) begin
              ways_0_metas_109_mru <= 1'b1;
            end
            if(_zz_112) begin
              ways_0_metas_110_mru <= 1'b1;
            end
            if(_zz_113) begin
              ways_0_metas_111_mru <= 1'b1;
            end
            if(_zz_114) begin
              ways_0_metas_112_mru <= 1'b1;
            end
            if(_zz_115) begin
              ways_0_metas_113_mru <= 1'b1;
            end
            if(_zz_116) begin
              ways_0_metas_114_mru <= 1'b1;
            end
            if(_zz_117) begin
              ways_0_metas_115_mru <= 1'b1;
            end
            if(_zz_118) begin
              ways_0_metas_116_mru <= 1'b1;
            end
            if(_zz_119) begin
              ways_0_metas_117_mru <= 1'b1;
            end
            if(_zz_120) begin
              ways_0_metas_118_mru <= 1'b1;
            end
            if(_zz_121) begin
              ways_0_metas_119_mru <= 1'b1;
            end
            if(_zz_122) begin
              ways_0_metas_120_mru <= 1'b1;
            end
            if(_zz_123) begin
              ways_0_metas_121_mru <= 1'b1;
            end
            if(_zz_124) begin
              ways_0_metas_122_mru <= 1'b1;
            end
            if(_zz_125) begin
              ways_0_metas_123_mru <= 1'b1;
            end
            if(_zz_126) begin
              ways_0_metas_124_mru <= 1'b1;
            end
            if(_zz_127) begin
              ways_0_metas_125_mru <= 1'b1;
            end
            if(_zz_128) begin
              ways_0_metas_126_mru <= 1'b1;
            end
            if(_zz_129) begin
              ways_0_metas_127_mru <= 1'b1;
            end
          end else begin
            if(when_ICache_l220) begin
              if(_zz_131) begin
                ways_0_metas_0_vld <= 1'b1;
              end
              if(_zz_132) begin
                ways_0_metas_1_vld <= 1'b1;
              end
              if(_zz_133) begin
                ways_0_metas_2_vld <= 1'b1;
              end
              if(_zz_134) begin
                ways_0_metas_3_vld <= 1'b1;
              end
              if(_zz_135) begin
                ways_0_metas_4_vld <= 1'b1;
              end
              if(_zz_136) begin
                ways_0_metas_5_vld <= 1'b1;
              end
              if(_zz_137) begin
                ways_0_metas_6_vld <= 1'b1;
              end
              if(_zz_138) begin
                ways_0_metas_7_vld <= 1'b1;
              end
              if(_zz_139) begin
                ways_0_metas_8_vld <= 1'b1;
              end
              if(_zz_140) begin
                ways_0_metas_9_vld <= 1'b1;
              end
              if(_zz_141) begin
                ways_0_metas_10_vld <= 1'b1;
              end
              if(_zz_142) begin
                ways_0_metas_11_vld <= 1'b1;
              end
              if(_zz_143) begin
                ways_0_metas_12_vld <= 1'b1;
              end
              if(_zz_144) begin
                ways_0_metas_13_vld <= 1'b1;
              end
              if(_zz_145) begin
                ways_0_metas_14_vld <= 1'b1;
              end
              if(_zz_146) begin
                ways_0_metas_15_vld <= 1'b1;
              end
              if(_zz_147) begin
                ways_0_metas_16_vld <= 1'b1;
              end
              if(_zz_148) begin
                ways_0_metas_17_vld <= 1'b1;
              end
              if(_zz_149) begin
                ways_0_metas_18_vld <= 1'b1;
              end
              if(_zz_150) begin
                ways_0_metas_19_vld <= 1'b1;
              end
              if(_zz_151) begin
                ways_0_metas_20_vld <= 1'b1;
              end
              if(_zz_152) begin
                ways_0_metas_21_vld <= 1'b1;
              end
              if(_zz_153) begin
                ways_0_metas_22_vld <= 1'b1;
              end
              if(_zz_154) begin
                ways_0_metas_23_vld <= 1'b1;
              end
              if(_zz_155) begin
                ways_0_metas_24_vld <= 1'b1;
              end
              if(_zz_156) begin
                ways_0_metas_25_vld <= 1'b1;
              end
              if(_zz_157) begin
                ways_0_metas_26_vld <= 1'b1;
              end
              if(_zz_158) begin
                ways_0_metas_27_vld <= 1'b1;
              end
              if(_zz_159) begin
                ways_0_metas_28_vld <= 1'b1;
              end
              if(_zz_160) begin
                ways_0_metas_29_vld <= 1'b1;
              end
              if(_zz_161) begin
                ways_0_metas_30_vld <= 1'b1;
              end
              if(_zz_162) begin
                ways_0_metas_31_vld <= 1'b1;
              end
              if(_zz_163) begin
                ways_0_metas_32_vld <= 1'b1;
              end
              if(_zz_164) begin
                ways_0_metas_33_vld <= 1'b1;
              end
              if(_zz_165) begin
                ways_0_metas_34_vld <= 1'b1;
              end
              if(_zz_166) begin
                ways_0_metas_35_vld <= 1'b1;
              end
              if(_zz_167) begin
                ways_0_metas_36_vld <= 1'b1;
              end
              if(_zz_168) begin
                ways_0_metas_37_vld <= 1'b1;
              end
              if(_zz_169) begin
                ways_0_metas_38_vld <= 1'b1;
              end
              if(_zz_170) begin
                ways_0_metas_39_vld <= 1'b1;
              end
              if(_zz_171) begin
                ways_0_metas_40_vld <= 1'b1;
              end
              if(_zz_172) begin
                ways_0_metas_41_vld <= 1'b1;
              end
              if(_zz_173) begin
                ways_0_metas_42_vld <= 1'b1;
              end
              if(_zz_174) begin
                ways_0_metas_43_vld <= 1'b1;
              end
              if(_zz_175) begin
                ways_0_metas_44_vld <= 1'b1;
              end
              if(_zz_176) begin
                ways_0_metas_45_vld <= 1'b1;
              end
              if(_zz_177) begin
                ways_0_metas_46_vld <= 1'b1;
              end
              if(_zz_178) begin
                ways_0_metas_47_vld <= 1'b1;
              end
              if(_zz_179) begin
                ways_0_metas_48_vld <= 1'b1;
              end
              if(_zz_180) begin
                ways_0_metas_49_vld <= 1'b1;
              end
              if(_zz_181) begin
                ways_0_metas_50_vld <= 1'b1;
              end
              if(_zz_182) begin
                ways_0_metas_51_vld <= 1'b1;
              end
              if(_zz_183) begin
                ways_0_metas_52_vld <= 1'b1;
              end
              if(_zz_184) begin
                ways_0_metas_53_vld <= 1'b1;
              end
              if(_zz_185) begin
                ways_0_metas_54_vld <= 1'b1;
              end
              if(_zz_186) begin
                ways_0_metas_55_vld <= 1'b1;
              end
              if(_zz_187) begin
                ways_0_metas_56_vld <= 1'b1;
              end
              if(_zz_188) begin
                ways_0_metas_57_vld <= 1'b1;
              end
              if(_zz_189) begin
                ways_0_metas_58_vld <= 1'b1;
              end
              if(_zz_190) begin
                ways_0_metas_59_vld <= 1'b1;
              end
              if(_zz_191) begin
                ways_0_metas_60_vld <= 1'b1;
              end
              if(_zz_192) begin
                ways_0_metas_61_vld <= 1'b1;
              end
              if(_zz_193) begin
                ways_0_metas_62_vld <= 1'b1;
              end
              if(_zz_194) begin
                ways_0_metas_63_vld <= 1'b1;
              end
              if(_zz_195) begin
                ways_0_metas_64_vld <= 1'b1;
              end
              if(_zz_196) begin
                ways_0_metas_65_vld <= 1'b1;
              end
              if(_zz_197) begin
                ways_0_metas_66_vld <= 1'b1;
              end
              if(_zz_198) begin
                ways_0_metas_67_vld <= 1'b1;
              end
              if(_zz_199) begin
                ways_0_metas_68_vld <= 1'b1;
              end
              if(_zz_200) begin
                ways_0_metas_69_vld <= 1'b1;
              end
              if(_zz_201) begin
                ways_0_metas_70_vld <= 1'b1;
              end
              if(_zz_202) begin
                ways_0_metas_71_vld <= 1'b1;
              end
              if(_zz_203) begin
                ways_0_metas_72_vld <= 1'b1;
              end
              if(_zz_204) begin
                ways_0_metas_73_vld <= 1'b1;
              end
              if(_zz_205) begin
                ways_0_metas_74_vld <= 1'b1;
              end
              if(_zz_206) begin
                ways_0_metas_75_vld <= 1'b1;
              end
              if(_zz_207) begin
                ways_0_metas_76_vld <= 1'b1;
              end
              if(_zz_208) begin
                ways_0_metas_77_vld <= 1'b1;
              end
              if(_zz_209) begin
                ways_0_metas_78_vld <= 1'b1;
              end
              if(_zz_210) begin
                ways_0_metas_79_vld <= 1'b1;
              end
              if(_zz_211) begin
                ways_0_metas_80_vld <= 1'b1;
              end
              if(_zz_212) begin
                ways_0_metas_81_vld <= 1'b1;
              end
              if(_zz_213) begin
                ways_0_metas_82_vld <= 1'b1;
              end
              if(_zz_214) begin
                ways_0_metas_83_vld <= 1'b1;
              end
              if(_zz_215) begin
                ways_0_metas_84_vld <= 1'b1;
              end
              if(_zz_216) begin
                ways_0_metas_85_vld <= 1'b1;
              end
              if(_zz_217) begin
                ways_0_metas_86_vld <= 1'b1;
              end
              if(_zz_218) begin
                ways_0_metas_87_vld <= 1'b1;
              end
              if(_zz_219) begin
                ways_0_metas_88_vld <= 1'b1;
              end
              if(_zz_220) begin
                ways_0_metas_89_vld <= 1'b1;
              end
              if(_zz_221) begin
                ways_0_metas_90_vld <= 1'b1;
              end
              if(_zz_222) begin
                ways_0_metas_91_vld <= 1'b1;
              end
              if(_zz_223) begin
                ways_0_metas_92_vld <= 1'b1;
              end
              if(_zz_224) begin
                ways_0_metas_93_vld <= 1'b1;
              end
              if(_zz_225) begin
                ways_0_metas_94_vld <= 1'b1;
              end
              if(_zz_226) begin
                ways_0_metas_95_vld <= 1'b1;
              end
              if(_zz_227) begin
                ways_0_metas_96_vld <= 1'b1;
              end
              if(_zz_228) begin
                ways_0_metas_97_vld <= 1'b1;
              end
              if(_zz_229) begin
                ways_0_metas_98_vld <= 1'b1;
              end
              if(_zz_230) begin
                ways_0_metas_99_vld <= 1'b1;
              end
              if(_zz_231) begin
                ways_0_metas_100_vld <= 1'b1;
              end
              if(_zz_232) begin
                ways_0_metas_101_vld <= 1'b1;
              end
              if(_zz_233) begin
                ways_0_metas_102_vld <= 1'b1;
              end
              if(_zz_234) begin
                ways_0_metas_103_vld <= 1'b1;
              end
              if(_zz_235) begin
                ways_0_metas_104_vld <= 1'b1;
              end
              if(_zz_236) begin
                ways_0_metas_105_vld <= 1'b1;
              end
              if(_zz_237) begin
                ways_0_metas_106_vld <= 1'b1;
              end
              if(_zz_238) begin
                ways_0_metas_107_vld <= 1'b1;
              end
              if(_zz_239) begin
                ways_0_metas_108_vld <= 1'b1;
              end
              if(_zz_240) begin
                ways_0_metas_109_vld <= 1'b1;
              end
              if(_zz_241) begin
                ways_0_metas_110_vld <= 1'b1;
              end
              if(_zz_242) begin
                ways_0_metas_111_vld <= 1'b1;
              end
              if(_zz_243) begin
                ways_0_metas_112_vld <= 1'b1;
              end
              if(_zz_244) begin
                ways_0_metas_113_vld <= 1'b1;
              end
              if(_zz_245) begin
                ways_0_metas_114_vld <= 1'b1;
              end
              if(_zz_246) begin
                ways_0_metas_115_vld <= 1'b1;
              end
              if(_zz_247) begin
                ways_0_metas_116_vld <= 1'b1;
              end
              if(_zz_248) begin
                ways_0_metas_117_vld <= 1'b1;
              end
              if(_zz_249) begin
                ways_0_metas_118_vld <= 1'b1;
              end
              if(_zz_250) begin
                ways_0_metas_119_vld <= 1'b1;
              end
              if(_zz_251) begin
                ways_0_metas_120_vld <= 1'b1;
              end
              if(_zz_252) begin
                ways_0_metas_121_vld <= 1'b1;
              end
              if(_zz_253) begin
                ways_0_metas_122_vld <= 1'b1;
              end
              if(_zz_254) begin
                ways_0_metas_123_vld <= 1'b1;
              end
              if(_zz_255) begin
                ways_0_metas_124_vld <= 1'b1;
              end
              if(_zz_256) begin
                ways_0_metas_125_vld <= 1'b1;
              end
              if(_zz_257) begin
                ways_0_metas_126_vld <= 1'b1;
              end
              if(_zz_258) begin
                ways_0_metas_127_vld <= 1'b1;
              end
            end
          end
        end
      end
      if(when_ICache_l225) begin
        if(_zz_131) begin
          ways_0_metas_0_tag <= cpu_tag_d1;
        end
        if(_zz_132) begin
          ways_0_metas_1_tag <= cpu_tag_d1;
        end
        if(_zz_133) begin
          ways_0_metas_2_tag <= cpu_tag_d1;
        end
        if(_zz_134) begin
          ways_0_metas_3_tag <= cpu_tag_d1;
        end
        if(_zz_135) begin
          ways_0_metas_4_tag <= cpu_tag_d1;
        end
        if(_zz_136) begin
          ways_0_metas_5_tag <= cpu_tag_d1;
        end
        if(_zz_137) begin
          ways_0_metas_6_tag <= cpu_tag_d1;
        end
        if(_zz_138) begin
          ways_0_metas_7_tag <= cpu_tag_d1;
        end
        if(_zz_139) begin
          ways_0_metas_8_tag <= cpu_tag_d1;
        end
        if(_zz_140) begin
          ways_0_metas_9_tag <= cpu_tag_d1;
        end
        if(_zz_141) begin
          ways_0_metas_10_tag <= cpu_tag_d1;
        end
        if(_zz_142) begin
          ways_0_metas_11_tag <= cpu_tag_d1;
        end
        if(_zz_143) begin
          ways_0_metas_12_tag <= cpu_tag_d1;
        end
        if(_zz_144) begin
          ways_0_metas_13_tag <= cpu_tag_d1;
        end
        if(_zz_145) begin
          ways_0_metas_14_tag <= cpu_tag_d1;
        end
        if(_zz_146) begin
          ways_0_metas_15_tag <= cpu_tag_d1;
        end
        if(_zz_147) begin
          ways_0_metas_16_tag <= cpu_tag_d1;
        end
        if(_zz_148) begin
          ways_0_metas_17_tag <= cpu_tag_d1;
        end
        if(_zz_149) begin
          ways_0_metas_18_tag <= cpu_tag_d1;
        end
        if(_zz_150) begin
          ways_0_metas_19_tag <= cpu_tag_d1;
        end
        if(_zz_151) begin
          ways_0_metas_20_tag <= cpu_tag_d1;
        end
        if(_zz_152) begin
          ways_0_metas_21_tag <= cpu_tag_d1;
        end
        if(_zz_153) begin
          ways_0_metas_22_tag <= cpu_tag_d1;
        end
        if(_zz_154) begin
          ways_0_metas_23_tag <= cpu_tag_d1;
        end
        if(_zz_155) begin
          ways_0_metas_24_tag <= cpu_tag_d1;
        end
        if(_zz_156) begin
          ways_0_metas_25_tag <= cpu_tag_d1;
        end
        if(_zz_157) begin
          ways_0_metas_26_tag <= cpu_tag_d1;
        end
        if(_zz_158) begin
          ways_0_metas_27_tag <= cpu_tag_d1;
        end
        if(_zz_159) begin
          ways_0_metas_28_tag <= cpu_tag_d1;
        end
        if(_zz_160) begin
          ways_0_metas_29_tag <= cpu_tag_d1;
        end
        if(_zz_161) begin
          ways_0_metas_30_tag <= cpu_tag_d1;
        end
        if(_zz_162) begin
          ways_0_metas_31_tag <= cpu_tag_d1;
        end
        if(_zz_163) begin
          ways_0_metas_32_tag <= cpu_tag_d1;
        end
        if(_zz_164) begin
          ways_0_metas_33_tag <= cpu_tag_d1;
        end
        if(_zz_165) begin
          ways_0_metas_34_tag <= cpu_tag_d1;
        end
        if(_zz_166) begin
          ways_0_metas_35_tag <= cpu_tag_d1;
        end
        if(_zz_167) begin
          ways_0_metas_36_tag <= cpu_tag_d1;
        end
        if(_zz_168) begin
          ways_0_metas_37_tag <= cpu_tag_d1;
        end
        if(_zz_169) begin
          ways_0_metas_38_tag <= cpu_tag_d1;
        end
        if(_zz_170) begin
          ways_0_metas_39_tag <= cpu_tag_d1;
        end
        if(_zz_171) begin
          ways_0_metas_40_tag <= cpu_tag_d1;
        end
        if(_zz_172) begin
          ways_0_metas_41_tag <= cpu_tag_d1;
        end
        if(_zz_173) begin
          ways_0_metas_42_tag <= cpu_tag_d1;
        end
        if(_zz_174) begin
          ways_0_metas_43_tag <= cpu_tag_d1;
        end
        if(_zz_175) begin
          ways_0_metas_44_tag <= cpu_tag_d1;
        end
        if(_zz_176) begin
          ways_0_metas_45_tag <= cpu_tag_d1;
        end
        if(_zz_177) begin
          ways_0_metas_46_tag <= cpu_tag_d1;
        end
        if(_zz_178) begin
          ways_0_metas_47_tag <= cpu_tag_d1;
        end
        if(_zz_179) begin
          ways_0_metas_48_tag <= cpu_tag_d1;
        end
        if(_zz_180) begin
          ways_0_metas_49_tag <= cpu_tag_d1;
        end
        if(_zz_181) begin
          ways_0_metas_50_tag <= cpu_tag_d1;
        end
        if(_zz_182) begin
          ways_0_metas_51_tag <= cpu_tag_d1;
        end
        if(_zz_183) begin
          ways_0_metas_52_tag <= cpu_tag_d1;
        end
        if(_zz_184) begin
          ways_0_metas_53_tag <= cpu_tag_d1;
        end
        if(_zz_185) begin
          ways_0_metas_54_tag <= cpu_tag_d1;
        end
        if(_zz_186) begin
          ways_0_metas_55_tag <= cpu_tag_d1;
        end
        if(_zz_187) begin
          ways_0_metas_56_tag <= cpu_tag_d1;
        end
        if(_zz_188) begin
          ways_0_metas_57_tag <= cpu_tag_d1;
        end
        if(_zz_189) begin
          ways_0_metas_58_tag <= cpu_tag_d1;
        end
        if(_zz_190) begin
          ways_0_metas_59_tag <= cpu_tag_d1;
        end
        if(_zz_191) begin
          ways_0_metas_60_tag <= cpu_tag_d1;
        end
        if(_zz_192) begin
          ways_0_metas_61_tag <= cpu_tag_d1;
        end
        if(_zz_193) begin
          ways_0_metas_62_tag <= cpu_tag_d1;
        end
        if(_zz_194) begin
          ways_0_metas_63_tag <= cpu_tag_d1;
        end
        if(_zz_195) begin
          ways_0_metas_64_tag <= cpu_tag_d1;
        end
        if(_zz_196) begin
          ways_0_metas_65_tag <= cpu_tag_d1;
        end
        if(_zz_197) begin
          ways_0_metas_66_tag <= cpu_tag_d1;
        end
        if(_zz_198) begin
          ways_0_metas_67_tag <= cpu_tag_d1;
        end
        if(_zz_199) begin
          ways_0_metas_68_tag <= cpu_tag_d1;
        end
        if(_zz_200) begin
          ways_0_metas_69_tag <= cpu_tag_d1;
        end
        if(_zz_201) begin
          ways_0_metas_70_tag <= cpu_tag_d1;
        end
        if(_zz_202) begin
          ways_0_metas_71_tag <= cpu_tag_d1;
        end
        if(_zz_203) begin
          ways_0_metas_72_tag <= cpu_tag_d1;
        end
        if(_zz_204) begin
          ways_0_metas_73_tag <= cpu_tag_d1;
        end
        if(_zz_205) begin
          ways_0_metas_74_tag <= cpu_tag_d1;
        end
        if(_zz_206) begin
          ways_0_metas_75_tag <= cpu_tag_d1;
        end
        if(_zz_207) begin
          ways_0_metas_76_tag <= cpu_tag_d1;
        end
        if(_zz_208) begin
          ways_0_metas_77_tag <= cpu_tag_d1;
        end
        if(_zz_209) begin
          ways_0_metas_78_tag <= cpu_tag_d1;
        end
        if(_zz_210) begin
          ways_0_metas_79_tag <= cpu_tag_d1;
        end
        if(_zz_211) begin
          ways_0_metas_80_tag <= cpu_tag_d1;
        end
        if(_zz_212) begin
          ways_0_metas_81_tag <= cpu_tag_d1;
        end
        if(_zz_213) begin
          ways_0_metas_82_tag <= cpu_tag_d1;
        end
        if(_zz_214) begin
          ways_0_metas_83_tag <= cpu_tag_d1;
        end
        if(_zz_215) begin
          ways_0_metas_84_tag <= cpu_tag_d1;
        end
        if(_zz_216) begin
          ways_0_metas_85_tag <= cpu_tag_d1;
        end
        if(_zz_217) begin
          ways_0_metas_86_tag <= cpu_tag_d1;
        end
        if(_zz_218) begin
          ways_0_metas_87_tag <= cpu_tag_d1;
        end
        if(_zz_219) begin
          ways_0_metas_88_tag <= cpu_tag_d1;
        end
        if(_zz_220) begin
          ways_0_metas_89_tag <= cpu_tag_d1;
        end
        if(_zz_221) begin
          ways_0_metas_90_tag <= cpu_tag_d1;
        end
        if(_zz_222) begin
          ways_0_metas_91_tag <= cpu_tag_d1;
        end
        if(_zz_223) begin
          ways_0_metas_92_tag <= cpu_tag_d1;
        end
        if(_zz_224) begin
          ways_0_metas_93_tag <= cpu_tag_d1;
        end
        if(_zz_225) begin
          ways_0_metas_94_tag <= cpu_tag_d1;
        end
        if(_zz_226) begin
          ways_0_metas_95_tag <= cpu_tag_d1;
        end
        if(_zz_227) begin
          ways_0_metas_96_tag <= cpu_tag_d1;
        end
        if(_zz_228) begin
          ways_0_metas_97_tag <= cpu_tag_d1;
        end
        if(_zz_229) begin
          ways_0_metas_98_tag <= cpu_tag_d1;
        end
        if(_zz_230) begin
          ways_0_metas_99_tag <= cpu_tag_d1;
        end
        if(_zz_231) begin
          ways_0_metas_100_tag <= cpu_tag_d1;
        end
        if(_zz_232) begin
          ways_0_metas_101_tag <= cpu_tag_d1;
        end
        if(_zz_233) begin
          ways_0_metas_102_tag <= cpu_tag_d1;
        end
        if(_zz_234) begin
          ways_0_metas_103_tag <= cpu_tag_d1;
        end
        if(_zz_235) begin
          ways_0_metas_104_tag <= cpu_tag_d1;
        end
        if(_zz_236) begin
          ways_0_metas_105_tag <= cpu_tag_d1;
        end
        if(_zz_237) begin
          ways_0_metas_106_tag <= cpu_tag_d1;
        end
        if(_zz_238) begin
          ways_0_metas_107_tag <= cpu_tag_d1;
        end
        if(_zz_239) begin
          ways_0_metas_108_tag <= cpu_tag_d1;
        end
        if(_zz_240) begin
          ways_0_metas_109_tag <= cpu_tag_d1;
        end
        if(_zz_241) begin
          ways_0_metas_110_tag <= cpu_tag_d1;
        end
        if(_zz_242) begin
          ways_0_metas_111_tag <= cpu_tag_d1;
        end
        if(_zz_243) begin
          ways_0_metas_112_tag <= cpu_tag_d1;
        end
        if(_zz_244) begin
          ways_0_metas_113_tag <= cpu_tag_d1;
        end
        if(_zz_245) begin
          ways_0_metas_114_tag <= cpu_tag_d1;
        end
        if(_zz_246) begin
          ways_0_metas_115_tag <= cpu_tag_d1;
        end
        if(_zz_247) begin
          ways_0_metas_116_tag <= cpu_tag_d1;
        end
        if(_zz_248) begin
          ways_0_metas_117_tag <= cpu_tag_d1;
        end
        if(_zz_249) begin
          ways_0_metas_118_tag <= cpu_tag_d1;
        end
        if(_zz_250) begin
          ways_0_metas_119_tag <= cpu_tag_d1;
        end
        if(_zz_251) begin
          ways_0_metas_120_tag <= cpu_tag_d1;
        end
        if(_zz_252) begin
          ways_0_metas_121_tag <= cpu_tag_d1;
        end
        if(_zz_253) begin
          ways_0_metas_122_tag <= cpu_tag_d1;
        end
        if(_zz_254) begin
          ways_0_metas_123_tag <= cpu_tag_d1;
        end
        if(_zz_255) begin
          ways_0_metas_124_tag <= cpu_tag_d1;
        end
        if(_zz_256) begin
          ways_0_metas_125_tag <= cpu_tag_d1;
        end
        if(_zz_257) begin
          ways_0_metas_126_tag <= cpu_tag_d1;
        end
        if(_zz_258) begin
          ways_0_metas_127_tag <= cpu_tag_d1;
        end
      end
      if(when_ICache_l230) begin
        cpu_cmd_ready_1 <= 1'b0;
      end else begin
        if(when_ICache_l233) begin
          cpu_cmd_ready_1 <= 1'b1;
        end
      end
      if(flush_busy) begin
        if(_zz_647) begin
          ways_1_metas_0_mru <= 1'b0;
        end
        if(_zz_648) begin
          ways_1_metas_1_mru <= 1'b0;
        end
        if(_zz_649) begin
          ways_1_metas_2_mru <= 1'b0;
        end
        if(_zz_650) begin
          ways_1_metas_3_mru <= 1'b0;
        end
        if(_zz_651) begin
          ways_1_metas_4_mru <= 1'b0;
        end
        if(_zz_652) begin
          ways_1_metas_5_mru <= 1'b0;
        end
        if(_zz_653) begin
          ways_1_metas_6_mru <= 1'b0;
        end
        if(_zz_654) begin
          ways_1_metas_7_mru <= 1'b0;
        end
        if(_zz_655) begin
          ways_1_metas_8_mru <= 1'b0;
        end
        if(_zz_656) begin
          ways_1_metas_9_mru <= 1'b0;
        end
        if(_zz_657) begin
          ways_1_metas_10_mru <= 1'b0;
        end
        if(_zz_658) begin
          ways_1_metas_11_mru <= 1'b0;
        end
        if(_zz_659) begin
          ways_1_metas_12_mru <= 1'b0;
        end
        if(_zz_660) begin
          ways_1_metas_13_mru <= 1'b0;
        end
        if(_zz_661) begin
          ways_1_metas_14_mru <= 1'b0;
        end
        if(_zz_662) begin
          ways_1_metas_15_mru <= 1'b0;
        end
        if(_zz_663) begin
          ways_1_metas_16_mru <= 1'b0;
        end
        if(_zz_664) begin
          ways_1_metas_17_mru <= 1'b0;
        end
        if(_zz_665) begin
          ways_1_metas_18_mru <= 1'b0;
        end
        if(_zz_666) begin
          ways_1_metas_19_mru <= 1'b0;
        end
        if(_zz_667) begin
          ways_1_metas_20_mru <= 1'b0;
        end
        if(_zz_668) begin
          ways_1_metas_21_mru <= 1'b0;
        end
        if(_zz_669) begin
          ways_1_metas_22_mru <= 1'b0;
        end
        if(_zz_670) begin
          ways_1_metas_23_mru <= 1'b0;
        end
        if(_zz_671) begin
          ways_1_metas_24_mru <= 1'b0;
        end
        if(_zz_672) begin
          ways_1_metas_25_mru <= 1'b0;
        end
        if(_zz_673) begin
          ways_1_metas_26_mru <= 1'b0;
        end
        if(_zz_674) begin
          ways_1_metas_27_mru <= 1'b0;
        end
        if(_zz_675) begin
          ways_1_metas_28_mru <= 1'b0;
        end
        if(_zz_676) begin
          ways_1_metas_29_mru <= 1'b0;
        end
        if(_zz_677) begin
          ways_1_metas_30_mru <= 1'b0;
        end
        if(_zz_678) begin
          ways_1_metas_31_mru <= 1'b0;
        end
        if(_zz_679) begin
          ways_1_metas_32_mru <= 1'b0;
        end
        if(_zz_680) begin
          ways_1_metas_33_mru <= 1'b0;
        end
        if(_zz_681) begin
          ways_1_metas_34_mru <= 1'b0;
        end
        if(_zz_682) begin
          ways_1_metas_35_mru <= 1'b0;
        end
        if(_zz_683) begin
          ways_1_metas_36_mru <= 1'b0;
        end
        if(_zz_684) begin
          ways_1_metas_37_mru <= 1'b0;
        end
        if(_zz_685) begin
          ways_1_metas_38_mru <= 1'b0;
        end
        if(_zz_686) begin
          ways_1_metas_39_mru <= 1'b0;
        end
        if(_zz_687) begin
          ways_1_metas_40_mru <= 1'b0;
        end
        if(_zz_688) begin
          ways_1_metas_41_mru <= 1'b0;
        end
        if(_zz_689) begin
          ways_1_metas_42_mru <= 1'b0;
        end
        if(_zz_690) begin
          ways_1_metas_43_mru <= 1'b0;
        end
        if(_zz_691) begin
          ways_1_metas_44_mru <= 1'b0;
        end
        if(_zz_692) begin
          ways_1_metas_45_mru <= 1'b0;
        end
        if(_zz_693) begin
          ways_1_metas_46_mru <= 1'b0;
        end
        if(_zz_694) begin
          ways_1_metas_47_mru <= 1'b0;
        end
        if(_zz_695) begin
          ways_1_metas_48_mru <= 1'b0;
        end
        if(_zz_696) begin
          ways_1_metas_49_mru <= 1'b0;
        end
        if(_zz_697) begin
          ways_1_metas_50_mru <= 1'b0;
        end
        if(_zz_698) begin
          ways_1_metas_51_mru <= 1'b0;
        end
        if(_zz_699) begin
          ways_1_metas_52_mru <= 1'b0;
        end
        if(_zz_700) begin
          ways_1_metas_53_mru <= 1'b0;
        end
        if(_zz_701) begin
          ways_1_metas_54_mru <= 1'b0;
        end
        if(_zz_702) begin
          ways_1_metas_55_mru <= 1'b0;
        end
        if(_zz_703) begin
          ways_1_metas_56_mru <= 1'b0;
        end
        if(_zz_704) begin
          ways_1_metas_57_mru <= 1'b0;
        end
        if(_zz_705) begin
          ways_1_metas_58_mru <= 1'b0;
        end
        if(_zz_706) begin
          ways_1_metas_59_mru <= 1'b0;
        end
        if(_zz_707) begin
          ways_1_metas_60_mru <= 1'b0;
        end
        if(_zz_708) begin
          ways_1_metas_61_mru <= 1'b0;
        end
        if(_zz_709) begin
          ways_1_metas_62_mru <= 1'b0;
        end
        if(_zz_710) begin
          ways_1_metas_63_mru <= 1'b0;
        end
        if(_zz_711) begin
          ways_1_metas_64_mru <= 1'b0;
        end
        if(_zz_712) begin
          ways_1_metas_65_mru <= 1'b0;
        end
        if(_zz_713) begin
          ways_1_metas_66_mru <= 1'b0;
        end
        if(_zz_714) begin
          ways_1_metas_67_mru <= 1'b0;
        end
        if(_zz_715) begin
          ways_1_metas_68_mru <= 1'b0;
        end
        if(_zz_716) begin
          ways_1_metas_69_mru <= 1'b0;
        end
        if(_zz_717) begin
          ways_1_metas_70_mru <= 1'b0;
        end
        if(_zz_718) begin
          ways_1_metas_71_mru <= 1'b0;
        end
        if(_zz_719) begin
          ways_1_metas_72_mru <= 1'b0;
        end
        if(_zz_720) begin
          ways_1_metas_73_mru <= 1'b0;
        end
        if(_zz_721) begin
          ways_1_metas_74_mru <= 1'b0;
        end
        if(_zz_722) begin
          ways_1_metas_75_mru <= 1'b0;
        end
        if(_zz_723) begin
          ways_1_metas_76_mru <= 1'b0;
        end
        if(_zz_724) begin
          ways_1_metas_77_mru <= 1'b0;
        end
        if(_zz_725) begin
          ways_1_metas_78_mru <= 1'b0;
        end
        if(_zz_726) begin
          ways_1_metas_79_mru <= 1'b0;
        end
        if(_zz_727) begin
          ways_1_metas_80_mru <= 1'b0;
        end
        if(_zz_728) begin
          ways_1_metas_81_mru <= 1'b0;
        end
        if(_zz_729) begin
          ways_1_metas_82_mru <= 1'b0;
        end
        if(_zz_730) begin
          ways_1_metas_83_mru <= 1'b0;
        end
        if(_zz_731) begin
          ways_1_metas_84_mru <= 1'b0;
        end
        if(_zz_732) begin
          ways_1_metas_85_mru <= 1'b0;
        end
        if(_zz_733) begin
          ways_1_metas_86_mru <= 1'b0;
        end
        if(_zz_734) begin
          ways_1_metas_87_mru <= 1'b0;
        end
        if(_zz_735) begin
          ways_1_metas_88_mru <= 1'b0;
        end
        if(_zz_736) begin
          ways_1_metas_89_mru <= 1'b0;
        end
        if(_zz_737) begin
          ways_1_metas_90_mru <= 1'b0;
        end
        if(_zz_738) begin
          ways_1_metas_91_mru <= 1'b0;
        end
        if(_zz_739) begin
          ways_1_metas_92_mru <= 1'b0;
        end
        if(_zz_740) begin
          ways_1_metas_93_mru <= 1'b0;
        end
        if(_zz_741) begin
          ways_1_metas_94_mru <= 1'b0;
        end
        if(_zz_742) begin
          ways_1_metas_95_mru <= 1'b0;
        end
        if(_zz_743) begin
          ways_1_metas_96_mru <= 1'b0;
        end
        if(_zz_744) begin
          ways_1_metas_97_mru <= 1'b0;
        end
        if(_zz_745) begin
          ways_1_metas_98_mru <= 1'b0;
        end
        if(_zz_746) begin
          ways_1_metas_99_mru <= 1'b0;
        end
        if(_zz_747) begin
          ways_1_metas_100_mru <= 1'b0;
        end
        if(_zz_748) begin
          ways_1_metas_101_mru <= 1'b0;
        end
        if(_zz_749) begin
          ways_1_metas_102_mru <= 1'b0;
        end
        if(_zz_750) begin
          ways_1_metas_103_mru <= 1'b0;
        end
        if(_zz_751) begin
          ways_1_metas_104_mru <= 1'b0;
        end
        if(_zz_752) begin
          ways_1_metas_105_mru <= 1'b0;
        end
        if(_zz_753) begin
          ways_1_metas_106_mru <= 1'b0;
        end
        if(_zz_754) begin
          ways_1_metas_107_mru <= 1'b0;
        end
        if(_zz_755) begin
          ways_1_metas_108_mru <= 1'b0;
        end
        if(_zz_756) begin
          ways_1_metas_109_mru <= 1'b0;
        end
        if(_zz_757) begin
          ways_1_metas_110_mru <= 1'b0;
        end
        if(_zz_758) begin
          ways_1_metas_111_mru <= 1'b0;
        end
        if(_zz_759) begin
          ways_1_metas_112_mru <= 1'b0;
        end
        if(_zz_760) begin
          ways_1_metas_113_mru <= 1'b0;
        end
        if(_zz_761) begin
          ways_1_metas_114_mru <= 1'b0;
        end
        if(_zz_762) begin
          ways_1_metas_115_mru <= 1'b0;
        end
        if(_zz_763) begin
          ways_1_metas_116_mru <= 1'b0;
        end
        if(_zz_764) begin
          ways_1_metas_117_mru <= 1'b0;
        end
        if(_zz_765) begin
          ways_1_metas_118_mru <= 1'b0;
        end
        if(_zz_766) begin
          ways_1_metas_119_mru <= 1'b0;
        end
        if(_zz_767) begin
          ways_1_metas_120_mru <= 1'b0;
        end
        if(_zz_768) begin
          ways_1_metas_121_mru <= 1'b0;
        end
        if(_zz_769) begin
          ways_1_metas_122_mru <= 1'b0;
        end
        if(_zz_770) begin
          ways_1_metas_123_mru <= 1'b0;
        end
        if(_zz_771) begin
          ways_1_metas_124_mru <= 1'b0;
        end
        if(_zz_772) begin
          ways_1_metas_125_mru <= 1'b0;
        end
        if(_zz_773) begin
          ways_1_metas_126_mru <= 1'b0;
        end
        if(_zz_774) begin
          ways_1_metas_127_mru <= 1'b0;
        end
        if(_zz_647) begin
          ways_1_metas_0_vld <= 1'b0;
        end
        if(_zz_648) begin
          ways_1_metas_1_vld <= 1'b0;
        end
        if(_zz_649) begin
          ways_1_metas_2_vld <= 1'b0;
        end
        if(_zz_650) begin
          ways_1_metas_3_vld <= 1'b0;
        end
        if(_zz_651) begin
          ways_1_metas_4_vld <= 1'b0;
        end
        if(_zz_652) begin
          ways_1_metas_5_vld <= 1'b0;
        end
        if(_zz_653) begin
          ways_1_metas_6_vld <= 1'b0;
        end
        if(_zz_654) begin
          ways_1_metas_7_vld <= 1'b0;
        end
        if(_zz_655) begin
          ways_1_metas_8_vld <= 1'b0;
        end
        if(_zz_656) begin
          ways_1_metas_9_vld <= 1'b0;
        end
        if(_zz_657) begin
          ways_1_metas_10_vld <= 1'b0;
        end
        if(_zz_658) begin
          ways_1_metas_11_vld <= 1'b0;
        end
        if(_zz_659) begin
          ways_1_metas_12_vld <= 1'b0;
        end
        if(_zz_660) begin
          ways_1_metas_13_vld <= 1'b0;
        end
        if(_zz_661) begin
          ways_1_metas_14_vld <= 1'b0;
        end
        if(_zz_662) begin
          ways_1_metas_15_vld <= 1'b0;
        end
        if(_zz_663) begin
          ways_1_metas_16_vld <= 1'b0;
        end
        if(_zz_664) begin
          ways_1_metas_17_vld <= 1'b0;
        end
        if(_zz_665) begin
          ways_1_metas_18_vld <= 1'b0;
        end
        if(_zz_666) begin
          ways_1_metas_19_vld <= 1'b0;
        end
        if(_zz_667) begin
          ways_1_metas_20_vld <= 1'b0;
        end
        if(_zz_668) begin
          ways_1_metas_21_vld <= 1'b0;
        end
        if(_zz_669) begin
          ways_1_metas_22_vld <= 1'b0;
        end
        if(_zz_670) begin
          ways_1_metas_23_vld <= 1'b0;
        end
        if(_zz_671) begin
          ways_1_metas_24_vld <= 1'b0;
        end
        if(_zz_672) begin
          ways_1_metas_25_vld <= 1'b0;
        end
        if(_zz_673) begin
          ways_1_metas_26_vld <= 1'b0;
        end
        if(_zz_674) begin
          ways_1_metas_27_vld <= 1'b0;
        end
        if(_zz_675) begin
          ways_1_metas_28_vld <= 1'b0;
        end
        if(_zz_676) begin
          ways_1_metas_29_vld <= 1'b0;
        end
        if(_zz_677) begin
          ways_1_metas_30_vld <= 1'b0;
        end
        if(_zz_678) begin
          ways_1_metas_31_vld <= 1'b0;
        end
        if(_zz_679) begin
          ways_1_metas_32_vld <= 1'b0;
        end
        if(_zz_680) begin
          ways_1_metas_33_vld <= 1'b0;
        end
        if(_zz_681) begin
          ways_1_metas_34_vld <= 1'b0;
        end
        if(_zz_682) begin
          ways_1_metas_35_vld <= 1'b0;
        end
        if(_zz_683) begin
          ways_1_metas_36_vld <= 1'b0;
        end
        if(_zz_684) begin
          ways_1_metas_37_vld <= 1'b0;
        end
        if(_zz_685) begin
          ways_1_metas_38_vld <= 1'b0;
        end
        if(_zz_686) begin
          ways_1_metas_39_vld <= 1'b0;
        end
        if(_zz_687) begin
          ways_1_metas_40_vld <= 1'b0;
        end
        if(_zz_688) begin
          ways_1_metas_41_vld <= 1'b0;
        end
        if(_zz_689) begin
          ways_1_metas_42_vld <= 1'b0;
        end
        if(_zz_690) begin
          ways_1_metas_43_vld <= 1'b0;
        end
        if(_zz_691) begin
          ways_1_metas_44_vld <= 1'b0;
        end
        if(_zz_692) begin
          ways_1_metas_45_vld <= 1'b0;
        end
        if(_zz_693) begin
          ways_1_metas_46_vld <= 1'b0;
        end
        if(_zz_694) begin
          ways_1_metas_47_vld <= 1'b0;
        end
        if(_zz_695) begin
          ways_1_metas_48_vld <= 1'b0;
        end
        if(_zz_696) begin
          ways_1_metas_49_vld <= 1'b0;
        end
        if(_zz_697) begin
          ways_1_metas_50_vld <= 1'b0;
        end
        if(_zz_698) begin
          ways_1_metas_51_vld <= 1'b0;
        end
        if(_zz_699) begin
          ways_1_metas_52_vld <= 1'b0;
        end
        if(_zz_700) begin
          ways_1_metas_53_vld <= 1'b0;
        end
        if(_zz_701) begin
          ways_1_metas_54_vld <= 1'b0;
        end
        if(_zz_702) begin
          ways_1_metas_55_vld <= 1'b0;
        end
        if(_zz_703) begin
          ways_1_metas_56_vld <= 1'b0;
        end
        if(_zz_704) begin
          ways_1_metas_57_vld <= 1'b0;
        end
        if(_zz_705) begin
          ways_1_metas_58_vld <= 1'b0;
        end
        if(_zz_706) begin
          ways_1_metas_59_vld <= 1'b0;
        end
        if(_zz_707) begin
          ways_1_metas_60_vld <= 1'b0;
        end
        if(_zz_708) begin
          ways_1_metas_61_vld <= 1'b0;
        end
        if(_zz_709) begin
          ways_1_metas_62_vld <= 1'b0;
        end
        if(_zz_710) begin
          ways_1_metas_63_vld <= 1'b0;
        end
        if(_zz_711) begin
          ways_1_metas_64_vld <= 1'b0;
        end
        if(_zz_712) begin
          ways_1_metas_65_vld <= 1'b0;
        end
        if(_zz_713) begin
          ways_1_metas_66_vld <= 1'b0;
        end
        if(_zz_714) begin
          ways_1_metas_67_vld <= 1'b0;
        end
        if(_zz_715) begin
          ways_1_metas_68_vld <= 1'b0;
        end
        if(_zz_716) begin
          ways_1_metas_69_vld <= 1'b0;
        end
        if(_zz_717) begin
          ways_1_metas_70_vld <= 1'b0;
        end
        if(_zz_718) begin
          ways_1_metas_71_vld <= 1'b0;
        end
        if(_zz_719) begin
          ways_1_metas_72_vld <= 1'b0;
        end
        if(_zz_720) begin
          ways_1_metas_73_vld <= 1'b0;
        end
        if(_zz_721) begin
          ways_1_metas_74_vld <= 1'b0;
        end
        if(_zz_722) begin
          ways_1_metas_75_vld <= 1'b0;
        end
        if(_zz_723) begin
          ways_1_metas_76_vld <= 1'b0;
        end
        if(_zz_724) begin
          ways_1_metas_77_vld <= 1'b0;
        end
        if(_zz_725) begin
          ways_1_metas_78_vld <= 1'b0;
        end
        if(_zz_726) begin
          ways_1_metas_79_vld <= 1'b0;
        end
        if(_zz_727) begin
          ways_1_metas_80_vld <= 1'b0;
        end
        if(_zz_728) begin
          ways_1_metas_81_vld <= 1'b0;
        end
        if(_zz_729) begin
          ways_1_metas_82_vld <= 1'b0;
        end
        if(_zz_730) begin
          ways_1_metas_83_vld <= 1'b0;
        end
        if(_zz_731) begin
          ways_1_metas_84_vld <= 1'b0;
        end
        if(_zz_732) begin
          ways_1_metas_85_vld <= 1'b0;
        end
        if(_zz_733) begin
          ways_1_metas_86_vld <= 1'b0;
        end
        if(_zz_734) begin
          ways_1_metas_87_vld <= 1'b0;
        end
        if(_zz_735) begin
          ways_1_metas_88_vld <= 1'b0;
        end
        if(_zz_736) begin
          ways_1_metas_89_vld <= 1'b0;
        end
        if(_zz_737) begin
          ways_1_metas_90_vld <= 1'b0;
        end
        if(_zz_738) begin
          ways_1_metas_91_vld <= 1'b0;
        end
        if(_zz_739) begin
          ways_1_metas_92_vld <= 1'b0;
        end
        if(_zz_740) begin
          ways_1_metas_93_vld <= 1'b0;
        end
        if(_zz_741) begin
          ways_1_metas_94_vld <= 1'b0;
        end
        if(_zz_742) begin
          ways_1_metas_95_vld <= 1'b0;
        end
        if(_zz_743) begin
          ways_1_metas_96_vld <= 1'b0;
        end
        if(_zz_744) begin
          ways_1_metas_97_vld <= 1'b0;
        end
        if(_zz_745) begin
          ways_1_metas_98_vld <= 1'b0;
        end
        if(_zz_746) begin
          ways_1_metas_99_vld <= 1'b0;
        end
        if(_zz_747) begin
          ways_1_metas_100_vld <= 1'b0;
        end
        if(_zz_748) begin
          ways_1_metas_101_vld <= 1'b0;
        end
        if(_zz_749) begin
          ways_1_metas_102_vld <= 1'b0;
        end
        if(_zz_750) begin
          ways_1_metas_103_vld <= 1'b0;
        end
        if(_zz_751) begin
          ways_1_metas_104_vld <= 1'b0;
        end
        if(_zz_752) begin
          ways_1_metas_105_vld <= 1'b0;
        end
        if(_zz_753) begin
          ways_1_metas_106_vld <= 1'b0;
        end
        if(_zz_754) begin
          ways_1_metas_107_vld <= 1'b0;
        end
        if(_zz_755) begin
          ways_1_metas_108_vld <= 1'b0;
        end
        if(_zz_756) begin
          ways_1_metas_109_vld <= 1'b0;
        end
        if(_zz_757) begin
          ways_1_metas_110_vld <= 1'b0;
        end
        if(_zz_758) begin
          ways_1_metas_111_vld <= 1'b0;
        end
        if(_zz_759) begin
          ways_1_metas_112_vld <= 1'b0;
        end
        if(_zz_760) begin
          ways_1_metas_113_vld <= 1'b0;
        end
        if(_zz_761) begin
          ways_1_metas_114_vld <= 1'b0;
        end
        if(_zz_762) begin
          ways_1_metas_115_vld <= 1'b0;
        end
        if(_zz_763) begin
          ways_1_metas_116_vld <= 1'b0;
        end
        if(_zz_764) begin
          ways_1_metas_117_vld <= 1'b0;
        end
        if(_zz_765) begin
          ways_1_metas_118_vld <= 1'b0;
        end
        if(_zz_766) begin
          ways_1_metas_119_vld <= 1'b0;
        end
        if(_zz_767) begin
          ways_1_metas_120_vld <= 1'b0;
        end
        if(_zz_768) begin
          ways_1_metas_121_vld <= 1'b0;
        end
        if(_zz_769) begin
          ways_1_metas_122_vld <= 1'b0;
        end
        if(_zz_770) begin
          ways_1_metas_123_vld <= 1'b0;
        end
        if(_zz_771) begin
          ways_1_metas_124_vld <= 1'b0;
        end
        if(_zz_772) begin
          ways_1_metas_125_vld <= 1'b0;
        end
        if(_zz_773) begin
          ways_1_metas_126_vld <= 1'b0;
        end
        if(_zz_774) begin
          ways_1_metas_127_vld <= 1'b0;
        end
      end else begin
        if(when_ICache_l210_1) begin
          if(cache_hit_1) begin
            if(_zz_389) begin
              ways_1_metas_0_mru <= 1'b1;
            end
            if(_zz_390) begin
              ways_1_metas_1_mru <= 1'b1;
            end
            if(_zz_391) begin
              ways_1_metas_2_mru <= 1'b1;
            end
            if(_zz_392) begin
              ways_1_metas_3_mru <= 1'b1;
            end
            if(_zz_393) begin
              ways_1_metas_4_mru <= 1'b1;
            end
            if(_zz_394) begin
              ways_1_metas_5_mru <= 1'b1;
            end
            if(_zz_395) begin
              ways_1_metas_6_mru <= 1'b1;
            end
            if(_zz_396) begin
              ways_1_metas_7_mru <= 1'b1;
            end
            if(_zz_397) begin
              ways_1_metas_8_mru <= 1'b1;
            end
            if(_zz_398) begin
              ways_1_metas_9_mru <= 1'b1;
            end
            if(_zz_399) begin
              ways_1_metas_10_mru <= 1'b1;
            end
            if(_zz_400) begin
              ways_1_metas_11_mru <= 1'b1;
            end
            if(_zz_401) begin
              ways_1_metas_12_mru <= 1'b1;
            end
            if(_zz_402) begin
              ways_1_metas_13_mru <= 1'b1;
            end
            if(_zz_403) begin
              ways_1_metas_14_mru <= 1'b1;
            end
            if(_zz_404) begin
              ways_1_metas_15_mru <= 1'b1;
            end
            if(_zz_405) begin
              ways_1_metas_16_mru <= 1'b1;
            end
            if(_zz_406) begin
              ways_1_metas_17_mru <= 1'b1;
            end
            if(_zz_407) begin
              ways_1_metas_18_mru <= 1'b1;
            end
            if(_zz_408) begin
              ways_1_metas_19_mru <= 1'b1;
            end
            if(_zz_409) begin
              ways_1_metas_20_mru <= 1'b1;
            end
            if(_zz_410) begin
              ways_1_metas_21_mru <= 1'b1;
            end
            if(_zz_411) begin
              ways_1_metas_22_mru <= 1'b1;
            end
            if(_zz_412) begin
              ways_1_metas_23_mru <= 1'b1;
            end
            if(_zz_413) begin
              ways_1_metas_24_mru <= 1'b1;
            end
            if(_zz_414) begin
              ways_1_metas_25_mru <= 1'b1;
            end
            if(_zz_415) begin
              ways_1_metas_26_mru <= 1'b1;
            end
            if(_zz_416) begin
              ways_1_metas_27_mru <= 1'b1;
            end
            if(_zz_417) begin
              ways_1_metas_28_mru <= 1'b1;
            end
            if(_zz_418) begin
              ways_1_metas_29_mru <= 1'b1;
            end
            if(_zz_419) begin
              ways_1_metas_30_mru <= 1'b1;
            end
            if(_zz_420) begin
              ways_1_metas_31_mru <= 1'b1;
            end
            if(_zz_421) begin
              ways_1_metas_32_mru <= 1'b1;
            end
            if(_zz_422) begin
              ways_1_metas_33_mru <= 1'b1;
            end
            if(_zz_423) begin
              ways_1_metas_34_mru <= 1'b1;
            end
            if(_zz_424) begin
              ways_1_metas_35_mru <= 1'b1;
            end
            if(_zz_425) begin
              ways_1_metas_36_mru <= 1'b1;
            end
            if(_zz_426) begin
              ways_1_metas_37_mru <= 1'b1;
            end
            if(_zz_427) begin
              ways_1_metas_38_mru <= 1'b1;
            end
            if(_zz_428) begin
              ways_1_metas_39_mru <= 1'b1;
            end
            if(_zz_429) begin
              ways_1_metas_40_mru <= 1'b1;
            end
            if(_zz_430) begin
              ways_1_metas_41_mru <= 1'b1;
            end
            if(_zz_431) begin
              ways_1_metas_42_mru <= 1'b1;
            end
            if(_zz_432) begin
              ways_1_metas_43_mru <= 1'b1;
            end
            if(_zz_433) begin
              ways_1_metas_44_mru <= 1'b1;
            end
            if(_zz_434) begin
              ways_1_metas_45_mru <= 1'b1;
            end
            if(_zz_435) begin
              ways_1_metas_46_mru <= 1'b1;
            end
            if(_zz_436) begin
              ways_1_metas_47_mru <= 1'b1;
            end
            if(_zz_437) begin
              ways_1_metas_48_mru <= 1'b1;
            end
            if(_zz_438) begin
              ways_1_metas_49_mru <= 1'b1;
            end
            if(_zz_439) begin
              ways_1_metas_50_mru <= 1'b1;
            end
            if(_zz_440) begin
              ways_1_metas_51_mru <= 1'b1;
            end
            if(_zz_441) begin
              ways_1_metas_52_mru <= 1'b1;
            end
            if(_zz_442) begin
              ways_1_metas_53_mru <= 1'b1;
            end
            if(_zz_443) begin
              ways_1_metas_54_mru <= 1'b1;
            end
            if(_zz_444) begin
              ways_1_metas_55_mru <= 1'b1;
            end
            if(_zz_445) begin
              ways_1_metas_56_mru <= 1'b1;
            end
            if(_zz_446) begin
              ways_1_metas_57_mru <= 1'b1;
            end
            if(_zz_447) begin
              ways_1_metas_58_mru <= 1'b1;
            end
            if(_zz_448) begin
              ways_1_metas_59_mru <= 1'b1;
            end
            if(_zz_449) begin
              ways_1_metas_60_mru <= 1'b1;
            end
            if(_zz_450) begin
              ways_1_metas_61_mru <= 1'b1;
            end
            if(_zz_451) begin
              ways_1_metas_62_mru <= 1'b1;
            end
            if(_zz_452) begin
              ways_1_metas_63_mru <= 1'b1;
            end
            if(_zz_453) begin
              ways_1_metas_64_mru <= 1'b1;
            end
            if(_zz_454) begin
              ways_1_metas_65_mru <= 1'b1;
            end
            if(_zz_455) begin
              ways_1_metas_66_mru <= 1'b1;
            end
            if(_zz_456) begin
              ways_1_metas_67_mru <= 1'b1;
            end
            if(_zz_457) begin
              ways_1_metas_68_mru <= 1'b1;
            end
            if(_zz_458) begin
              ways_1_metas_69_mru <= 1'b1;
            end
            if(_zz_459) begin
              ways_1_metas_70_mru <= 1'b1;
            end
            if(_zz_460) begin
              ways_1_metas_71_mru <= 1'b1;
            end
            if(_zz_461) begin
              ways_1_metas_72_mru <= 1'b1;
            end
            if(_zz_462) begin
              ways_1_metas_73_mru <= 1'b1;
            end
            if(_zz_463) begin
              ways_1_metas_74_mru <= 1'b1;
            end
            if(_zz_464) begin
              ways_1_metas_75_mru <= 1'b1;
            end
            if(_zz_465) begin
              ways_1_metas_76_mru <= 1'b1;
            end
            if(_zz_466) begin
              ways_1_metas_77_mru <= 1'b1;
            end
            if(_zz_467) begin
              ways_1_metas_78_mru <= 1'b1;
            end
            if(_zz_468) begin
              ways_1_metas_79_mru <= 1'b1;
            end
            if(_zz_469) begin
              ways_1_metas_80_mru <= 1'b1;
            end
            if(_zz_470) begin
              ways_1_metas_81_mru <= 1'b1;
            end
            if(_zz_471) begin
              ways_1_metas_82_mru <= 1'b1;
            end
            if(_zz_472) begin
              ways_1_metas_83_mru <= 1'b1;
            end
            if(_zz_473) begin
              ways_1_metas_84_mru <= 1'b1;
            end
            if(_zz_474) begin
              ways_1_metas_85_mru <= 1'b1;
            end
            if(_zz_475) begin
              ways_1_metas_86_mru <= 1'b1;
            end
            if(_zz_476) begin
              ways_1_metas_87_mru <= 1'b1;
            end
            if(_zz_477) begin
              ways_1_metas_88_mru <= 1'b1;
            end
            if(_zz_478) begin
              ways_1_metas_89_mru <= 1'b1;
            end
            if(_zz_479) begin
              ways_1_metas_90_mru <= 1'b1;
            end
            if(_zz_480) begin
              ways_1_metas_91_mru <= 1'b1;
            end
            if(_zz_481) begin
              ways_1_metas_92_mru <= 1'b1;
            end
            if(_zz_482) begin
              ways_1_metas_93_mru <= 1'b1;
            end
            if(_zz_483) begin
              ways_1_metas_94_mru <= 1'b1;
            end
            if(_zz_484) begin
              ways_1_metas_95_mru <= 1'b1;
            end
            if(_zz_485) begin
              ways_1_metas_96_mru <= 1'b1;
            end
            if(_zz_486) begin
              ways_1_metas_97_mru <= 1'b1;
            end
            if(_zz_487) begin
              ways_1_metas_98_mru <= 1'b1;
            end
            if(_zz_488) begin
              ways_1_metas_99_mru <= 1'b1;
            end
            if(_zz_489) begin
              ways_1_metas_100_mru <= 1'b1;
            end
            if(_zz_490) begin
              ways_1_metas_101_mru <= 1'b1;
            end
            if(_zz_491) begin
              ways_1_metas_102_mru <= 1'b1;
            end
            if(_zz_492) begin
              ways_1_metas_103_mru <= 1'b1;
            end
            if(_zz_493) begin
              ways_1_metas_104_mru <= 1'b1;
            end
            if(_zz_494) begin
              ways_1_metas_105_mru <= 1'b1;
            end
            if(_zz_495) begin
              ways_1_metas_106_mru <= 1'b1;
            end
            if(_zz_496) begin
              ways_1_metas_107_mru <= 1'b1;
            end
            if(_zz_497) begin
              ways_1_metas_108_mru <= 1'b1;
            end
            if(_zz_498) begin
              ways_1_metas_109_mru <= 1'b1;
            end
            if(_zz_499) begin
              ways_1_metas_110_mru <= 1'b1;
            end
            if(_zz_500) begin
              ways_1_metas_111_mru <= 1'b1;
            end
            if(_zz_501) begin
              ways_1_metas_112_mru <= 1'b1;
            end
            if(_zz_502) begin
              ways_1_metas_113_mru <= 1'b1;
            end
            if(_zz_503) begin
              ways_1_metas_114_mru <= 1'b1;
            end
            if(_zz_504) begin
              ways_1_metas_115_mru <= 1'b1;
            end
            if(_zz_505) begin
              ways_1_metas_116_mru <= 1'b1;
            end
            if(_zz_506) begin
              ways_1_metas_117_mru <= 1'b1;
            end
            if(_zz_507) begin
              ways_1_metas_118_mru <= 1'b1;
            end
            if(_zz_508) begin
              ways_1_metas_119_mru <= 1'b1;
            end
            if(_zz_509) begin
              ways_1_metas_120_mru <= 1'b1;
            end
            if(_zz_510) begin
              ways_1_metas_121_mru <= 1'b1;
            end
            if(_zz_511) begin
              ways_1_metas_122_mru <= 1'b1;
            end
            if(_zz_512) begin
              ways_1_metas_123_mru <= 1'b1;
            end
            if(_zz_513) begin
              ways_1_metas_124_mru <= 1'b1;
            end
            if(_zz_514) begin
              ways_1_metas_125_mru <= 1'b1;
            end
            if(_zz_515) begin
              ways_1_metas_126_mru <= 1'b1;
            end
            if(_zz_516) begin
              ways_1_metas_127_mru <= 1'b1;
            end
          end else begin
            if(_zz_389) begin
              ways_1_metas_0_mru <= 1'b0;
            end
            if(_zz_390) begin
              ways_1_metas_1_mru <= 1'b0;
            end
            if(_zz_391) begin
              ways_1_metas_2_mru <= 1'b0;
            end
            if(_zz_392) begin
              ways_1_metas_3_mru <= 1'b0;
            end
            if(_zz_393) begin
              ways_1_metas_4_mru <= 1'b0;
            end
            if(_zz_394) begin
              ways_1_metas_5_mru <= 1'b0;
            end
            if(_zz_395) begin
              ways_1_metas_6_mru <= 1'b0;
            end
            if(_zz_396) begin
              ways_1_metas_7_mru <= 1'b0;
            end
            if(_zz_397) begin
              ways_1_metas_8_mru <= 1'b0;
            end
            if(_zz_398) begin
              ways_1_metas_9_mru <= 1'b0;
            end
            if(_zz_399) begin
              ways_1_metas_10_mru <= 1'b0;
            end
            if(_zz_400) begin
              ways_1_metas_11_mru <= 1'b0;
            end
            if(_zz_401) begin
              ways_1_metas_12_mru <= 1'b0;
            end
            if(_zz_402) begin
              ways_1_metas_13_mru <= 1'b0;
            end
            if(_zz_403) begin
              ways_1_metas_14_mru <= 1'b0;
            end
            if(_zz_404) begin
              ways_1_metas_15_mru <= 1'b0;
            end
            if(_zz_405) begin
              ways_1_metas_16_mru <= 1'b0;
            end
            if(_zz_406) begin
              ways_1_metas_17_mru <= 1'b0;
            end
            if(_zz_407) begin
              ways_1_metas_18_mru <= 1'b0;
            end
            if(_zz_408) begin
              ways_1_metas_19_mru <= 1'b0;
            end
            if(_zz_409) begin
              ways_1_metas_20_mru <= 1'b0;
            end
            if(_zz_410) begin
              ways_1_metas_21_mru <= 1'b0;
            end
            if(_zz_411) begin
              ways_1_metas_22_mru <= 1'b0;
            end
            if(_zz_412) begin
              ways_1_metas_23_mru <= 1'b0;
            end
            if(_zz_413) begin
              ways_1_metas_24_mru <= 1'b0;
            end
            if(_zz_414) begin
              ways_1_metas_25_mru <= 1'b0;
            end
            if(_zz_415) begin
              ways_1_metas_26_mru <= 1'b0;
            end
            if(_zz_416) begin
              ways_1_metas_27_mru <= 1'b0;
            end
            if(_zz_417) begin
              ways_1_metas_28_mru <= 1'b0;
            end
            if(_zz_418) begin
              ways_1_metas_29_mru <= 1'b0;
            end
            if(_zz_419) begin
              ways_1_metas_30_mru <= 1'b0;
            end
            if(_zz_420) begin
              ways_1_metas_31_mru <= 1'b0;
            end
            if(_zz_421) begin
              ways_1_metas_32_mru <= 1'b0;
            end
            if(_zz_422) begin
              ways_1_metas_33_mru <= 1'b0;
            end
            if(_zz_423) begin
              ways_1_metas_34_mru <= 1'b0;
            end
            if(_zz_424) begin
              ways_1_metas_35_mru <= 1'b0;
            end
            if(_zz_425) begin
              ways_1_metas_36_mru <= 1'b0;
            end
            if(_zz_426) begin
              ways_1_metas_37_mru <= 1'b0;
            end
            if(_zz_427) begin
              ways_1_metas_38_mru <= 1'b0;
            end
            if(_zz_428) begin
              ways_1_metas_39_mru <= 1'b0;
            end
            if(_zz_429) begin
              ways_1_metas_40_mru <= 1'b0;
            end
            if(_zz_430) begin
              ways_1_metas_41_mru <= 1'b0;
            end
            if(_zz_431) begin
              ways_1_metas_42_mru <= 1'b0;
            end
            if(_zz_432) begin
              ways_1_metas_43_mru <= 1'b0;
            end
            if(_zz_433) begin
              ways_1_metas_44_mru <= 1'b0;
            end
            if(_zz_434) begin
              ways_1_metas_45_mru <= 1'b0;
            end
            if(_zz_435) begin
              ways_1_metas_46_mru <= 1'b0;
            end
            if(_zz_436) begin
              ways_1_metas_47_mru <= 1'b0;
            end
            if(_zz_437) begin
              ways_1_metas_48_mru <= 1'b0;
            end
            if(_zz_438) begin
              ways_1_metas_49_mru <= 1'b0;
            end
            if(_zz_439) begin
              ways_1_metas_50_mru <= 1'b0;
            end
            if(_zz_440) begin
              ways_1_metas_51_mru <= 1'b0;
            end
            if(_zz_441) begin
              ways_1_metas_52_mru <= 1'b0;
            end
            if(_zz_442) begin
              ways_1_metas_53_mru <= 1'b0;
            end
            if(_zz_443) begin
              ways_1_metas_54_mru <= 1'b0;
            end
            if(_zz_444) begin
              ways_1_metas_55_mru <= 1'b0;
            end
            if(_zz_445) begin
              ways_1_metas_56_mru <= 1'b0;
            end
            if(_zz_446) begin
              ways_1_metas_57_mru <= 1'b0;
            end
            if(_zz_447) begin
              ways_1_metas_58_mru <= 1'b0;
            end
            if(_zz_448) begin
              ways_1_metas_59_mru <= 1'b0;
            end
            if(_zz_449) begin
              ways_1_metas_60_mru <= 1'b0;
            end
            if(_zz_450) begin
              ways_1_metas_61_mru <= 1'b0;
            end
            if(_zz_451) begin
              ways_1_metas_62_mru <= 1'b0;
            end
            if(_zz_452) begin
              ways_1_metas_63_mru <= 1'b0;
            end
            if(_zz_453) begin
              ways_1_metas_64_mru <= 1'b0;
            end
            if(_zz_454) begin
              ways_1_metas_65_mru <= 1'b0;
            end
            if(_zz_455) begin
              ways_1_metas_66_mru <= 1'b0;
            end
            if(_zz_456) begin
              ways_1_metas_67_mru <= 1'b0;
            end
            if(_zz_457) begin
              ways_1_metas_68_mru <= 1'b0;
            end
            if(_zz_458) begin
              ways_1_metas_69_mru <= 1'b0;
            end
            if(_zz_459) begin
              ways_1_metas_70_mru <= 1'b0;
            end
            if(_zz_460) begin
              ways_1_metas_71_mru <= 1'b0;
            end
            if(_zz_461) begin
              ways_1_metas_72_mru <= 1'b0;
            end
            if(_zz_462) begin
              ways_1_metas_73_mru <= 1'b0;
            end
            if(_zz_463) begin
              ways_1_metas_74_mru <= 1'b0;
            end
            if(_zz_464) begin
              ways_1_metas_75_mru <= 1'b0;
            end
            if(_zz_465) begin
              ways_1_metas_76_mru <= 1'b0;
            end
            if(_zz_466) begin
              ways_1_metas_77_mru <= 1'b0;
            end
            if(_zz_467) begin
              ways_1_metas_78_mru <= 1'b0;
            end
            if(_zz_468) begin
              ways_1_metas_79_mru <= 1'b0;
            end
            if(_zz_469) begin
              ways_1_metas_80_mru <= 1'b0;
            end
            if(_zz_470) begin
              ways_1_metas_81_mru <= 1'b0;
            end
            if(_zz_471) begin
              ways_1_metas_82_mru <= 1'b0;
            end
            if(_zz_472) begin
              ways_1_metas_83_mru <= 1'b0;
            end
            if(_zz_473) begin
              ways_1_metas_84_mru <= 1'b0;
            end
            if(_zz_474) begin
              ways_1_metas_85_mru <= 1'b0;
            end
            if(_zz_475) begin
              ways_1_metas_86_mru <= 1'b0;
            end
            if(_zz_476) begin
              ways_1_metas_87_mru <= 1'b0;
            end
            if(_zz_477) begin
              ways_1_metas_88_mru <= 1'b0;
            end
            if(_zz_478) begin
              ways_1_metas_89_mru <= 1'b0;
            end
            if(_zz_479) begin
              ways_1_metas_90_mru <= 1'b0;
            end
            if(_zz_480) begin
              ways_1_metas_91_mru <= 1'b0;
            end
            if(_zz_481) begin
              ways_1_metas_92_mru <= 1'b0;
            end
            if(_zz_482) begin
              ways_1_metas_93_mru <= 1'b0;
            end
            if(_zz_483) begin
              ways_1_metas_94_mru <= 1'b0;
            end
            if(_zz_484) begin
              ways_1_metas_95_mru <= 1'b0;
            end
            if(_zz_485) begin
              ways_1_metas_96_mru <= 1'b0;
            end
            if(_zz_486) begin
              ways_1_metas_97_mru <= 1'b0;
            end
            if(_zz_487) begin
              ways_1_metas_98_mru <= 1'b0;
            end
            if(_zz_488) begin
              ways_1_metas_99_mru <= 1'b0;
            end
            if(_zz_489) begin
              ways_1_metas_100_mru <= 1'b0;
            end
            if(_zz_490) begin
              ways_1_metas_101_mru <= 1'b0;
            end
            if(_zz_491) begin
              ways_1_metas_102_mru <= 1'b0;
            end
            if(_zz_492) begin
              ways_1_metas_103_mru <= 1'b0;
            end
            if(_zz_493) begin
              ways_1_metas_104_mru <= 1'b0;
            end
            if(_zz_494) begin
              ways_1_metas_105_mru <= 1'b0;
            end
            if(_zz_495) begin
              ways_1_metas_106_mru <= 1'b0;
            end
            if(_zz_496) begin
              ways_1_metas_107_mru <= 1'b0;
            end
            if(_zz_497) begin
              ways_1_metas_108_mru <= 1'b0;
            end
            if(_zz_498) begin
              ways_1_metas_109_mru <= 1'b0;
            end
            if(_zz_499) begin
              ways_1_metas_110_mru <= 1'b0;
            end
            if(_zz_500) begin
              ways_1_metas_111_mru <= 1'b0;
            end
            if(_zz_501) begin
              ways_1_metas_112_mru <= 1'b0;
            end
            if(_zz_502) begin
              ways_1_metas_113_mru <= 1'b0;
            end
            if(_zz_503) begin
              ways_1_metas_114_mru <= 1'b0;
            end
            if(_zz_504) begin
              ways_1_metas_115_mru <= 1'b0;
            end
            if(_zz_505) begin
              ways_1_metas_116_mru <= 1'b0;
            end
            if(_zz_506) begin
              ways_1_metas_117_mru <= 1'b0;
            end
            if(_zz_507) begin
              ways_1_metas_118_mru <= 1'b0;
            end
            if(_zz_508) begin
              ways_1_metas_119_mru <= 1'b0;
            end
            if(_zz_509) begin
              ways_1_metas_120_mru <= 1'b0;
            end
            if(_zz_510) begin
              ways_1_metas_121_mru <= 1'b0;
            end
            if(_zz_511) begin
              ways_1_metas_122_mru <= 1'b0;
            end
            if(_zz_512) begin
              ways_1_metas_123_mru <= 1'b0;
            end
            if(_zz_513) begin
              ways_1_metas_124_mru <= 1'b0;
            end
            if(_zz_514) begin
              ways_1_metas_125_mru <= 1'b0;
            end
            if(_zz_515) begin
              ways_1_metas_126_mru <= 1'b0;
            end
            if(_zz_516) begin
              ways_1_metas_127_mru <= 1'b0;
            end
          end
        end else begin
          if(when_ICache_l217_1) begin
            if(_zz_389) begin
              ways_1_metas_0_mru <= 1'b1;
            end
            if(_zz_390) begin
              ways_1_metas_1_mru <= 1'b1;
            end
            if(_zz_391) begin
              ways_1_metas_2_mru <= 1'b1;
            end
            if(_zz_392) begin
              ways_1_metas_3_mru <= 1'b1;
            end
            if(_zz_393) begin
              ways_1_metas_4_mru <= 1'b1;
            end
            if(_zz_394) begin
              ways_1_metas_5_mru <= 1'b1;
            end
            if(_zz_395) begin
              ways_1_metas_6_mru <= 1'b1;
            end
            if(_zz_396) begin
              ways_1_metas_7_mru <= 1'b1;
            end
            if(_zz_397) begin
              ways_1_metas_8_mru <= 1'b1;
            end
            if(_zz_398) begin
              ways_1_metas_9_mru <= 1'b1;
            end
            if(_zz_399) begin
              ways_1_metas_10_mru <= 1'b1;
            end
            if(_zz_400) begin
              ways_1_metas_11_mru <= 1'b1;
            end
            if(_zz_401) begin
              ways_1_metas_12_mru <= 1'b1;
            end
            if(_zz_402) begin
              ways_1_metas_13_mru <= 1'b1;
            end
            if(_zz_403) begin
              ways_1_metas_14_mru <= 1'b1;
            end
            if(_zz_404) begin
              ways_1_metas_15_mru <= 1'b1;
            end
            if(_zz_405) begin
              ways_1_metas_16_mru <= 1'b1;
            end
            if(_zz_406) begin
              ways_1_metas_17_mru <= 1'b1;
            end
            if(_zz_407) begin
              ways_1_metas_18_mru <= 1'b1;
            end
            if(_zz_408) begin
              ways_1_metas_19_mru <= 1'b1;
            end
            if(_zz_409) begin
              ways_1_metas_20_mru <= 1'b1;
            end
            if(_zz_410) begin
              ways_1_metas_21_mru <= 1'b1;
            end
            if(_zz_411) begin
              ways_1_metas_22_mru <= 1'b1;
            end
            if(_zz_412) begin
              ways_1_metas_23_mru <= 1'b1;
            end
            if(_zz_413) begin
              ways_1_metas_24_mru <= 1'b1;
            end
            if(_zz_414) begin
              ways_1_metas_25_mru <= 1'b1;
            end
            if(_zz_415) begin
              ways_1_metas_26_mru <= 1'b1;
            end
            if(_zz_416) begin
              ways_1_metas_27_mru <= 1'b1;
            end
            if(_zz_417) begin
              ways_1_metas_28_mru <= 1'b1;
            end
            if(_zz_418) begin
              ways_1_metas_29_mru <= 1'b1;
            end
            if(_zz_419) begin
              ways_1_metas_30_mru <= 1'b1;
            end
            if(_zz_420) begin
              ways_1_metas_31_mru <= 1'b1;
            end
            if(_zz_421) begin
              ways_1_metas_32_mru <= 1'b1;
            end
            if(_zz_422) begin
              ways_1_metas_33_mru <= 1'b1;
            end
            if(_zz_423) begin
              ways_1_metas_34_mru <= 1'b1;
            end
            if(_zz_424) begin
              ways_1_metas_35_mru <= 1'b1;
            end
            if(_zz_425) begin
              ways_1_metas_36_mru <= 1'b1;
            end
            if(_zz_426) begin
              ways_1_metas_37_mru <= 1'b1;
            end
            if(_zz_427) begin
              ways_1_metas_38_mru <= 1'b1;
            end
            if(_zz_428) begin
              ways_1_metas_39_mru <= 1'b1;
            end
            if(_zz_429) begin
              ways_1_metas_40_mru <= 1'b1;
            end
            if(_zz_430) begin
              ways_1_metas_41_mru <= 1'b1;
            end
            if(_zz_431) begin
              ways_1_metas_42_mru <= 1'b1;
            end
            if(_zz_432) begin
              ways_1_metas_43_mru <= 1'b1;
            end
            if(_zz_433) begin
              ways_1_metas_44_mru <= 1'b1;
            end
            if(_zz_434) begin
              ways_1_metas_45_mru <= 1'b1;
            end
            if(_zz_435) begin
              ways_1_metas_46_mru <= 1'b1;
            end
            if(_zz_436) begin
              ways_1_metas_47_mru <= 1'b1;
            end
            if(_zz_437) begin
              ways_1_metas_48_mru <= 1'b1;
            end
            if(_zz_438) begin
              ways_1_metas_49_mru <= 1'b1;
            end
            if(_zz_439) begin
              ways_1_metas_50_mru <= 1'b1;
            end
            if(_zz_440) begin
              ways_1_metas_51_mru <= 1'b1;
            end
            if(_zz_441) begin
              ways_1_metas_52_mru <= 1'b1;
            end
            if(_zz_442) begin
              ways_1_metas_53_mru <= 1'b1;
            end
            if(_zz_443) begin
              ways_1_metas_54_mru <= 1'b1;
            end
            if(_zz_444) begin
              ways_1_metas_55_mru <= 1'b1;
            end
            if(_zz_445) begin
              ways_1_metas_56_mru <= 1'b1;
            end
            if(_zz_446) begin
              ways_1_metas_57_mru <= 1'b1;
            end
            if(_zz_447) begin
              ways_1_metas_58_mru <= 1'b1;
            end
            if(_zz_448) begin
              ways_1_metas_59_mru <= 1'b1;
            end
            if(_zz_449) begin
              ways_1_metas_60_mru <= 1'b1;
            end
            if(_zz_450) begin
              ways_1_metas_61_mru <= 1'b1;
            end
            if(_zz_451) begin
              ways_1_metas_62_mru <= 1'b1;
            end
            if(_zz_452) begin
              ways_1_metas_63_mru <= 1'b1;
            end
            if(_zz_453) begin
              ways_1_metas_64_mru <= 1'b1;
            end
            if(_zz_454) begin
              ways_1_metas_65_mru <= 1'b1;
            end
            if(_zz_455) begin
              ways_1_metas_66_mru <= 1'b1;
            end
            if(_zz_456) begin
              ways_1_metas_67_mru <= 1'b1;
            end
            if(_zz_457) begin
              ways_1_metas_68_mru <= 1'b1;
            end
            if(_zz_458) begin
              ways_1_metas_69_mru <= 1'b1;
            end
            if(_zz_459) begin
              ways_1_metas_70_mru <= 1'b1;
            end
            if(_zz_460) begin
              ways_1_metas_71_mru <= 1'b1;
            end
            if(_zz_461) begin
              ways_1_metas_72_mru <= 1'b1;
            end
            if(_zz_462) begin
              ways_1_metas_73_mru <= 1'b1;
            end
            if(_zz_463) begin
              ways_1_metas_74_mru <= 1'b1;
            end
            if(_zz_464) begin
              ways_1_metas_75_mru <= 1'b1;
            end
            if(_zz_465) begin
              ways_1_metas_76_mru <= 1'b1;
            end
            if(_zz_466) begin
              ways_1_metas_77_mru <= 1'b1;
            end
            if(_zz_467) begin
              ways_1_metas_78_mru <= 1'b1;
            end
            if(_zz_468) begin
              ways_1_metas_79_mru <= 1'b1;
            end
            if(_zz_469) begin
              ways_1_metas_80_mru <= 1'b1;
            end
            if(_zz_470) begin
              ways_1_metas_81_mru <= 1'b1;
            end
            if(_zz_471) begin
              ways_1_metas_82_mru <= 1'b1;
            end
            if(_zz_472) begin
              ways_1_metas_83_mru <= 1'b1;
            end
            if(_zz_473) begin
              ways_1_metas_84_mru <= 1'b1;
            end
            if(_zz_474) begin
              ways_1_metas_85_mru <= 1'b1;
            end
            if(_zz_475) begin
              ways_1_metas_86_mru <= 1'b1;
            end
            if(_zz_476) begin
              ways_1_metas_87_mru <= 1'b1;
            end
            if(_zz_477) begin
              ways_1_metas_88_mru <= 1'b1;
            end
            if(_zz_478) begin
              ways_1_metas_89_mru <= 1'b1;
            end
            if(_zz_479) begin
              ways_1_metas_90_mru <= 1'b1;
            end
            if(_zz_480) begin
              ways_1_metas_91_mru <= 1'b1;
            end
            if(_zz_481) begin
              ways_1_metas_92_mru <= 1'b1;
            end
            if(_zz_482) begin
              ways_1_metas_93_mru <= 1'b1;
            end
            if(_zz_483) begin
              ways_1_metas_94_mru <= 1'b1;
            end
            if(_zz_484) begin
              ways_1_metas_95_mru <= 1'b1;
            end
            if(_zz_485) begin
              ways_1_metas_96_mru <= 1'b1;
            end
            if(_zz_486) begin
              ways_1_metas_97_mru <= 1'b1;
            end
            if(_zz_487) begin
              ways_1_metas_98_mru <= 1'b1;
            end
            if(_zz_488) begin
              ways_1_metas_99_mru <= 1'b1;
            end
            if(_zz_489) begin
              ways_1_metas_100_mru <= 1'b1;
            end
            if(_zz_490) begin
              ways_1_metas_101_mru <= 1'b1;
            end
            if(_zz_491) begin
              ways_1_metas_102_mru <= 1'b1;
            end
            if(_zz_492) begin
              ways_1_metas_103_mru <= 1'b1;
            end
            if(_zz_493) begin
              ways_1_metas_104_mru <= 1'b1;
            end
            if(_zz_494) begin
              ways_1_metas_105_mru <= 1'b1;
            end
            if(_zz_495) begin
              ways_1_metas_106_mru <= 1'b1;
            end
            if(_zz_496) begin
              ways_1_metas_107_mru <= 1'b1;
            end
            if(_zz_497) begin
              ways_1_metas_108_mru <= 1'b1;
            end
            if(_zz_498) begin
              ways_1_metas_109_mru <= 1'b1;
            end
            if(_zz_499) begin
              ways_1_metas_110_mru <= 1'b1;
            end
            if(_zz_500) begin
              ways_1_metas_111_mru <= 1'b1;
            end
            if(_zz_501) begin
              ways_1_metas_112_mru <= 1'b1;
            end
            if(_zz_502) begin
              ways_1_metas_113_mru <= 1'b1;
            end
            if(_zz_503) begin
              ways_1_metas_114_mru <= 1'b1;
            end
            if(_zz_504) begin
              ways_1_metas_115_mru <= 1'b1;
            end
            if(_zz_505) begin
              ways_1_metas_116_mru <= 1'b1;
            end
            if(_zz_506) begin
              ways_1_metas_117_mru <= 1'b1;
            end
            if(_zz_507) begin
              ways_1_metas_118_mru <= 1'b1;
            end
            if(_zz_508) begin
              ways_1_metas_119_mru <= 1'b1;
            end
            if(_zz_509) begin
              ways_1_metas_120_mru <= 1'b1;
            end
            if(_zz_510) begin
              ways_1_metas_121_mru <= 1'b1;
            end
            if(_zz_511) begin
              ways_1_metas_122_mru <= 1'b1;
            end
            if(_zz_512) begin
              ways_1_metas_123_mru <= 1'b1;
            end
            if(_zz_513) begin
              ways_1_metas_124_mru <= 1'b1;
            end
            if(_zz_514) begin
              ways_1_metas_125_mru <= 1'b1;
            end
            if(_zz_515) begin
              ways_1_metas_126_mru <= 1'b1;
            end
            if(_zz_516) begin
              ways_1_metas_127_mru <= 1'b1;
            end
          end else begin
            if(when_ICache_l220_1) begin
              if(_zz_518) begin
                ways_1_metas_0_vld <= 1'b1;
              end
              if(_zz_519) begin
                ways_1_metas_1_vld <= 1'b1;
              end
              if(_zz_520) begin
                ways_1_metas_2_vld <= 1'b1;
              end
              if(_zz_521) begin
                ways_1_metas_3_vld <= 1'b1;
              end
              if(_zz_522) begin
                ways_1_metas_4_vld <= 1'b1;
              end
              if(_zz_523) begin
                ways_1_metas_5_vld <= 1'b1;
              end
              if(_zz_524) begin
                ways_1_metas_6_vld <= 1'b1;
              end
              if(_zz_525) begin
                ways_1_metas_7_vld <= 1'b1;
              end
              if(_zz_526) begin
                ways_1_metas_8_vld <= 1'b1;
              end
              if(_zz_527) begin
                ways_1_metas_9_vld <= 1'b1;
              end
              if(_zz_528) begin
                ways_1_metas_10_vld <= 1'b1;
              end
              if(_zz_529) begin
                ways_1_metas_11_vld <= 1'b1;
              end
              if(_zz_530) begin
                ways_1_metas_12_vld <= 1'b1;
              end
              if(_zz_531) begin
                ways_1_metas_13_vld <= 1'b1;
              end
              if(_zz_532) begin
                ways_1_metas_14_vld <= 1'b1;
              end
              if(_zz_533) begin
                ways_1_metas_15_vld <= 1'b1;
              end
              if(_zz_534) begin
                ways_1_metas_16_vld <= 1'b1;
              end
              if(_zz_535) begin
                ways_1_metas_17_vld <= 1'b1;
              end
              if(_zz_536) begin
                ways_1_metas_18_vld <= 1'b1;
              end
              if(_zz_537) begin
                ways_1_metas_19_vld <= 1'b1;
              end
              if(_zz_538) begin
                ways_1_metas_20_vld <= 1'b1;
              end
              if(_zz_539) begin
                ways_1_metas_21_vld <= 1'b1;
              end
              if(_zz_540) begin
                ways_1_metas_22_vld <= 1'b1;
              end
              if(_zz_541) begin
                ways_1_metas_23_vld <= 1'b1;
              end
              if(_zz_542) begin
                ways_1_metas_24_vld <= 1'b1;
              end
              if(_zz_543) begin
                ways_1_metas_25_vld <= 1'b1;
              end
              if(_zz_544) begin
                ways_1_metas_26_vld <= 1'b1;
              end
              if(_zz_545) begin
                ways_1_metas_27_vld <= 1'b1;
              end
              if(_zz_546) begin
                ways_1_metas_28_vld <= 1'b1;
              end
              if(_zz_547) begin
                ways_1_metas_29_vld <= 1'b1;
              end
              if(_zz_548) begin
                ways_1_metas_30_vld <= 1'b1;
              end
              if(_zz_549) begin
                ways_1_metas_31_vld <= 1'b1;
              end
              if(_zz_550) begin
                ways_1_metas_32_vld <= 1'b1;
              end
              if(_zz_551) begin
                ways_1_metas_33_vld <= 1'b1;
              end
              if(_zz_552) begin
                ways_1_metas_34_vld <= 1'b1;
              end
              if(_zz_553) begin
                ways_1_metas_35_vld <= 1'b1;
              end
              if(_zz_554) begin
                ways_1_metas_36_vld <= 1'b1;
              end
              if(_zz_555) begin
                ways_1_metas_37_vld <= 1'b1;
              end
              if(_zz_556) begin
                ways_1_metas_38_vld <= 1'b1;
              end
              if(_zz_557) begin
                ways_1_metas_39_vld <= 1'b1;
              end
              if(_zz_558) begin
                ways_1_metas_40_vld <= 1'b1;
              end
              if(_zz_559) begin
                ways_1_metas_41_vld <= 1'b1;
              end
              if(_zz_560) begin
                ways_1_metas_42_vld <= 1'b1;
              end
              if(_zz_561) begin
                ways_1_metas_43_vld <= 1'b1;
              end
              if(_zz_562) begin
                ways_1_metas_44_vld <= 1'b1;
              end
              if(_zz_563) begin
                ways_1_metas_45_vld <= 1'b1;
              end
              if(_zz_564) begin
                ways_1_metas_46_vld <= 1'b1;
              end
              if(_zz_565) begin
                ways_1_metas_47_vld <= 1'b1;
              end
              if(_zz_566) begin
                ways_1_metas_48_vld <= 1'b1;
              end
              if(_zz_567) begin
                ways_1_metas_49_vld <= 1'b1;
              end
              if(_zz_568) begin
                ways_1_metas_50_vld <= 1'b1;
              end
              if(_zz_569) begin
                ways_1_metas_51_vld <= 1'b1;
              end
              if(_zz_570) begin
                ways_1_metas_52_vld <= 1'b1;
              end
              if(_zz_571) begin
                ways_1_metas_53_vld <= 1'b1;
              end
              if(_zz_572) begin
                ways_1_metas_54_vld <= 1'b1;
              end
              if(_zz_573) begin
                ways_1_metas_55_vld <= 1'b1;
              end
              if(_zz_574) begin
                ways_1_metas_56_vld <= 1'b1;
              end
              if(_zz_575) begin
                ways_1_metas_57_vld <= 1'b1;
              end
              if(_zz_576) begin
                ways_1_metas_58_vld <= 1'b1;
              end
              if(_zz_577) begin
                ways_1_metas_59_vld <= 1'b1;
              end
              if(_zz_578) begin
                ways_1_metas_60_vld <= 1'b1;
              end
              if(_zz_579) begin
                ways_1_metas_61_vld <= 1'b1;
              end
              if(_zz_580) begin
                ways_1_metas_62_vld <= 1'b1;
              end
              if(_zz_581) begin
                ways_1_metas_63_vld <= 1'b1;
              end
              if(_zz_582) begin
                ways_1_metas_64_vld <= 1'b1;
              end
              if(_zz_583) begin
                ways_1_metas_65_vld <= 1'b1;
              end
              if(_zz_584) begin
                ways_1_metas_66_vld <= 1'b1;
              end
              if(_zz_585) begin
                ways_1_metas_67_vld <= 1'b1;
              end
              if(_zz_586) begin
                ways_1_metas_68_vld <= 1'b1;
              end
              if(_zz_587) begin
                ways_1_metas_69_vld <= 1'b1;
              end
              if(_zz_588) begin
                ways_1_metas_70_vld <= 1'b1;
              end
              if(_zz_589) begin
                ways_1_metas_71_vld <= 1'b1;
              end
              if(_zz_590) begin
                ways_1_metas_72_vld <= 1'b1;
              end
              if(_zz_591) begin
                ways_1_metas_73_vld <= 1'b1;
              end
              if(_zz_592) begin
                ways_1_metas_74_vld <= 1'b1;
              end
              if(_zz_593) begin
                ways_1_metas_75_vld <= 1'b1;
              end
              if(_zz_594) begin
                ways_1_metas_76_vld <= 1'b1;
              end
              if(_zz_595) begin
                ways_1_metas_77_vld <= 1'b1;
              end
              if(_zz_596) begin
                ways_1_metas_78_vld <= 1'b1;
              end
              if(_zz_597) begin
                ways_1_metas_79_vld <= 1'b1;
              end
              if(_zz_598) begin
                ways_1_metas_80_vld <= 1'b1;
              end
              if(_zz_599) begin
                ways_1_metas_81_vld <= 1'b1;
              end
              if(_zz_600) begin
                ways_1_metas_82_vld <= 1'b1;
              end
              if(_zz_601) begin
                ways_1_metas_83_vld <= 1'b1;
              end
              if(_zz_602) begin
                ways_1_metas_84_vld <= 1'b1;
              end
              if(_zz_603) begin
                ways_1_metas_85_vld <= 1'b1;
              end
              if(_zz_604) begin
                ways_1_metas_86_vld <= 1'b1;
              end
              if(_zz_605) begin
                ways_1_metas_87_vld <= 1'b1;
              end
              if(_zz_606) begin
                ways_1_metas_88_vld <= 1'b1;
              end
              if(_zz_607) begin
                ways_1_metas_89_vld <= 1'b1;
              end
              if(_zz_608) begin
                ways_1_metas_90_vld <= 1'b1;
              end
              if(_zz_609) begin
                ways_1_metas_91_vld <= 1'b1;
              end
              if(_zz_610) begin
                ways_1_metas_92_vld <= 1'b1;
              end
              if(_zz_611) begin
                ways_1_metas_93_vld <= 1'b1;
              end
              if(_zz_612) begin
                ways_1_metas_94_vld <= 1'b1;
              end
              if(_zz_613) begin
                ways_1_metas_95_vld <= 1'b1;
              end
              if(_zz_614) begin
                ways_1_metas_96_vld <= 1'b1;
              end
              if(_zz_615) begin
                ways_1_metas_97_vld <= 1'b1;
              end
              if(_zz_616) begin
                ways_1_metas_98_vld <= 1'b1;
              end
              if(_zz_617) begin
                ways_1_metas_99_vld <= 1'b1;
              end
              if(_zz_618) begin
                ways_1_metas_100_vld <= 1'b1;
              end
              if(_zz_619) begin
                ways_1_metas_101_vld <= 1'b1;
              end
              if(_zz_620) begin
                ways_1_metas_102_vld <= 1'b1;
              end
              if(_zz_621) begin
                ways_1_metas_103_vld <= 1'b1;
              end
              if(_zz_622) begin
                ways_1_metas_104_vld <= 1'b1;
              end
              if(_zz_623) begin
                ways_1_metas_105_vld <= 1'b1;
              end
              if(_zz_624) begin
                ways_1_metas_106_vld <= 1'b1;
              end
              if(_zz_625) begin
                ways_1_metas_107_vld <= 1'b1;
              end
              if(_zz_626) begin
                ways_1_metas_108_vld <= 1'b1;
              end
              if(_zz_627) begin
                ways_1_metas_109_vld <= 1'b1;
              end
              if(_zz_628) begin
                ways_1_metas_110_vld <= 1'b1;
              end
              if(_zz_629) begin
                ways_1_metas_111_vld <= 1'b1;
              end
              if(_zz_630) begin
                ways_1_metas_112_vld <= 1'b1;
              end
              if(_zz_631) begin
                ways_1_metas_113_vld <= 1'b1;
              end
              if(_zz_632) begin
                ways_1_metas_114_vld <= 1'b1;
              end
              if(_zz_633) begin
                ways_1_metas_115_vld <= 1'b1;
              end
              if(_zz_634) begin
                ways_1_metas_116_vld <= 1'b1;
              end
              if(_zz_635) begin
                ways_1_metas_117_vld <= 1'b1;
              end
              if(_zz_636) begin
                ways_1_metas_118_vld <= 1'b1;
              end
              if(_zz_637) begin
                ways_1_metas_119_vld <= 1'b1;
              end
              if(_zz_638) begin
                ways_1_metas_120_vld <= 1'b1;
              end
              if(_zz_639) begin
                ways_1_metas_121_vld <= 1'b1;
              end
              if(_zz_640) begin
                ways_1_metas_122_vld <= 1'b1;
              end
              if(_zz_641) begin
                ways_1_metas_123_vld <= 1'b1;
              end
              if(_zz_642) begin
                ways_1_metas_124_vld <= 1'b1;
              end
              if(_zz_643) begin
                ways_1_metas_125_vld <= 1'b1;
              end
              if(_zz_644) begin
                ways_1_metas_126_vld <= 1'b1;
              end
              if(_zz_645) begin
                ways_1_metas_127_vld <= 1'b1;
              end
            end
          end
        end
      end
      if(when_ICache_l225_1) begin
        if(_zz_518) begin
          ways_1_metas_0_tag <= cpu_tag_d1;
        end
        if(_zz_519) begin
          ways_1_metas_1_tag <= cpu_tag_d1;
        end
        if(_zz_520) begin
          ways_1_metas_2_tag <= cpu_tag_d1;
        end
        if(_zz_521) begin
          ways_1_metas_3_tag <= cpu_tag_d1;
        end
        if(_zz_522) begin
          ways_1_metas_4_tag <= cpu_tag_d1;
        end
        if(_zz_523) begin
          ways_1_metas_5_tag <= cpu_tag_d1;
        end
        if(_zz_524) begin
          ways_1_metas_6_tag <= cpu_tag_d1;
        end
        if(_zz_525) begin
          ways_1_metas_7_tag <= cpu_tag_d1;
        end
        if(_zz_526) begin
          ways_1_metas_8_tag <= cpu_tag_d1;
        end
        if(_zz_527) begin
          ways_1_metas_9_tag <= cpu_tag_d1;
        end
        if(_zz_528) begin
          ways_1_metas_10_tag <= cpu_tag_d1;
        end
        if(_zz_529) begin
          ways_1_metas_11_tag <= cpu_tag_d1;
        end
        if(_zz_530) begin
          ways_1_metas_12_tag <= cpu_tag_d1;
        end
        if(_zz_531) begin
          ways_1_metas_13_tag <= cpu_tag_d1;
        end
        if(_zz_532) begin
          ways_1_metas_14_tag <= cpu_tag_d1;
        end
        if(_zz_533) begin
          ways_1_metas_15_tag <= cpu_tag_d1;
        end
        if(_zz_534) begin
          ways_1_metas_16_tag <= cpu_tag_d1;
        end
        if(_zz_535) begin
          ways_1_metas_17_tag <= cpu_tag_d1;
        end
        if(_zz_536) begin
          ways_1_metas_18_tag <= cpu_tag_d1;
        end
        if(_zz_537) begin
          ways_1_metas_19_tag <= cpu_tag_d1;
        end
        if(_zz_538) begin
          ways_1_metas_20_tag <= cpu_tag_d1;
        end
        if(_zz_539) begin
          ways_1_metas_21_tag <= cpu_tag_d1;
        end
        if(_zz_540) begin
          ways_1_metas_22_tag <= cpu_tag_d1;
        end
        if(_zz_541) begin
          ways_1_metas_23_tag <= cpu_tag_d1;
        end
        if(_zz_542) begin
          ways_1_metas_24_tag <= cpu_tag_d1;
        end
        if(_zz_543) begin
          ways_1_metas_25_tag <= cpu_tag_d1;
        end
        if(_zz_544) begin
          ways_1_metas_26_tag <= cpu_tag_d1;
        end
        if(_zz_545) begin
          ways_1_metas_27_tag <= cpu_tag_d1;
        end
        if(_zz_546) begin
          ways_1_metas_28_tag <= cpu_tag_d1;
        end
        if(_zz_547) begin
          ways_1_metas_29_tag <= cpu_tag_d1;
        end
        if(_zz_548) begin
          ways_1_metas_30_tag <= cpu_tag_d1;
        end
        if(_zz_549) begin
          ways_1_metas_31_tag <= cpu_tag_d1;
        end
        if(_zz_550) begin
          ways_1_metas_32_tag <= cpu_tag_d1;
        end
        if(_zz_551) begin
          ways_1_metas_33_tag <= cpu_tag_d1;
        end
        if(_zz_552) begin
          ways_1_metas_34_tag <= cpu_tag_d1;
        end
        if(_zz_553) begin
          ways_1_metas_35_tag <= cpu_tag_d1;
        end
        if(_zz_554) begin
          ways_1_metas_36_tag <= cpu_tag_d1;
        end
        if(_zz_555) begin
          ways_1_metas_37_tag <= cpu_tag_d1;
        end
        if(_zz_556) begin
          ways_1_metas_38_tag <= cpu_tag_d1;
        end
        if(_zz_557) begin
          ways_1_metas_39_tag <= cpu_tag_d1;
        end
        if(_zz_558) begin
          ways_1_metas_40_tag <= cpu_tag_d1;
        end
        if(_zz_559) begin
          ways_1_metas_41_tag <= cpu_tag_d1;
        end
        if(_zz_560) begin
          ways_1_metas_42_tag <= cpu_tag_d1;
        end
        if(_zz_561) begin
          ways_1_metas_43_tag <= cpu_tag_d1;
        end
        if(_zz_562) begin
          ways_1_metas_44_tag <= cpu_tag_d1;
        end
        if(_zz_563) begin
          ways_1_metas_45_tag <= cpu_tag_d1;
        end
        if(_zz_564) begin
          ways_1_metas_46_tag <= cpu_tag_d1;
        end
        if(_zz_565) begin
          ways_1_metas_47_tag <= cpu_tag_d1;
        end
        if(_zz_566) begin
          ways_1_metas_48_tag <= cpu_tag_d1;
        end
        if(_zz_567) begin
          ways_1_metas_49_tag <= cpu_tag_d1;
        end
        if(_zz_568) begin
          ways_1_metas_50_tag <= cpu_tag_d1;
        end
        if(_zz_569) begin
          ways_1_metas_51_tag <= cpu_tag_d1;
        end
        if(_zz_570) begin
          ways_1_metas_52_tag <= cpu_tag_d1;
        end
        if(_zz_571) begin
          ways_1_metas_53_tag <= cpu_tag_d1;
        end
        if(_zz_572) begin
          ways_1_metas_54_tag <= cpu_tag_d1;
        end
        if(_zz_573) begin
          ways_1_metas_55_tag <= cpu_tag_d1;
        end
        if(_zz_574) begin
          ways_1_metas_56_tag <= cpu_tag_d1;
        end
        if(_zz_575) begin
          ways_1_metas_57_tag <= cpu_tag_d1;
        end
        if(_zz_576) begin
          ways_1_metas_58_tag <= cpu_tag_d1;
        end
        if(_zz_577) begin
          ways_1_metas_59_tag <= cpu_tag_d1;
        end
        if(_zz_578) begin
          ways_1_metas_60_tag <= cpu_tag_d1;
        end
        if(_zz_579) begin
          ways_1_metas_61_tag <= cpu_tag_d1;
        end
        if(_zz_580) begin
          ways_1_metas_62_tag <= cpu_tag_d1;
        end
        if(_zz_581) begin
          ways_1_metas_63_tag <= cpu_tag_d1;
        end
        if(_zz_582) begin
          ways_1_metas_64_tag <= cpu_tag_d1;
        end
        if(_zz_583) begin
          ways_1_metas_65_tag <= cpu_tag_d1;
        end
        if(_zz_584) begin
          ways_1_metas_66_tag <= cpu_tag_d1;
        end
        if(_zz_585) begin
          ways_1_metas_67_tag <= cpu_tag_d1;
        end
        if(_zz_586) begin
          ways_1_metas_68_tag <= cpu_tag_d1;
        end
        if(_zz_587) begin
          ways_1_metas_69_tag <= cpu_tag_d1;
        end
        if(_zz_588) begin
          ways_1_metas_70_tag <= cpu_tag_d1;
        end
        if(_zz_589) begin
          ways_1_metas_71_tag <= cpu_tag_d1;
        end
        if(_zz_590) begin
          ways_1_metas_72_tag <= cpu_tag_d1;
        end
        if(_zz_591) begin
          ways_1_metas_73_tag <= cpu_tag_d1;
        end
        if(_zz_592) begin
          ways_1_metas_74_tag <= cpu_tag_d1;
        end
        if(_zz_593) begin
          ways_1_metas_75_tag <= cpu_tag_d1;
        end
        if(_zz_594) begin
          ways_1_metas_76_tag <= cpu_tag_d1;
        end
        if(_zz_595) begin
          ways_1_metas_77_tag <= cpu_tag_d1;
        end
        if(_zz_596) begin
          ways_1_metas_78_tag <= cpu_tag_d1;
        end
        if(_zz_597) begin
          ways_1_metas_79_tag <= cpu_tag_d1;
        end
        if(_zz_598) begin
          ways_1_metas_80_tag <= cpu_tag_d1;
        end
        if(_zz_599) begin
          ways_1_metas_81_tag <= cpu_tag_d1;
        end
        if(_zz_600) begin
          ways_1_metas_82_tag <= cpu_tag_d1;
        end
        if(_zz_601) begin
          ways_1_metas_83_tag <= cpu_tag_d1;
        end
        if(_zz_602) begin
          ways_1_metas_84_tag <= cpu_tag_d1;
        end
        if(_zz_603) begin
          ways_1_metas_85_tag <= cpu_tag_d1;
        end
        if(_zz_604) begin
          ways_1_metas_86_tag <= cpu_tag_d1;
        end
        if(_zz_605) begin
          ways_1_metas_87_tag <= cpu_tag_d1;
        end
        if(_zz_606) begin
          ways_1_metas_88_tag <= cpu_tag_d1;
        end
        if(_zz_607) begin
          ways_1_metas_89_tag <= cpu_tag_d1;
        end
        if(_zz_608) begin
          ways_1_metas_90_tag <= cpu_tag_d1;
        end
        if(_zz_609) begin
          ways_1_metas_91_tag <= cpu_tag_d1;
        end
        if(_zz_610) begin
          ways_1_metas_92_tag <= cpu_tag_d1;
        end
        if(_zz_611) begin
          ways_1_metas_93_tag <= cpu_tag_d1;
        end
        if(_zz_612) begin
          ways_1_metas_94_tag <= cpu_tag_d1;
        end
        if(_zz_613) begin
          ways_1_metas_95_tag <= cpu_tag_d1;
        end
        if(_zz_614) begin
          ways_1_metas_96_tag <= cpu_tag_d1;
        end
        if(_zz_615) begin
          ways_1_metas_97_tag <= cpu_tag_d1;
        end
        if(_zz_616) begin
          ways_1_metas_98_tag <= cpu_tag_d1;
        end
        if(_zz_617) begin
          ways_1_metas_99_tag <= cpu_tag_d1;
        end
        if(_zz_618) begin
          ways_1_metas_100_tag <= cpu_tag_d1;
        end
        if(_zz_619) begin
          ways_1_metas_101_tag <= cpu_tag_d1;
        end
        if(_zz_620) begin
          ways_1_metas_102_tag <= cpu_tag_d1;
        end
        if(_zz_621) begin
          ways_1_metas_103_tag <= cpu_tag_d1;
        end
        if(_zz_622) begin
          ways_1_metas_104_tag <= cpu_tag_d1;
        end
        if(_zz_623) begin
          ways_1_metas_105_tag <= cpu_tag_d1;
        end
        if(_zz_624) begin
          ways_1_metas_106_tag <= cpu_tag_d1;
        end
        if(_zz_625) begin
          ways_1_metas_107_tag <= cpu_tag_d1;
        end
        if(_zz_626) begin
          ways_1_metas_108_tag <= cpu_tag_d1;
        end
        if(_zz_627) begin
          ways_1_metas_109_tag <= cpu_tag_d1;
        end
        if(_zz_628) begin
          ways_1_metas_110_tag <= cpu_tag_d1;
        end
        if(_zz_629) begin
          ways_1_metas_111_tag <= cpu_tag_d1;
        end
        if(_zz_630) begin
          ways_1_metas_112_tag <= cpu_tag_d1;
        end
        if(_zz_631) begin
          ways_1_metas_113_tag <= cpu_tag_d1;
        end
        if(_zz_632) begin
          ways_1_metas_114_tag <= cpu_tag_d1;
        end
        if(_zz_633) begin
          ways_1_metas_115_tag <= cpu_tag_d1;
        end
        if(_zz_634) begin
          ways_1_metas_116_tag <= cpu_tag_d1;
        end
        if(_zz_635) begin
          ways_1_metas_117_tag <= cpu_tag_d1;
        end
        if(_zz_636) begin
          ways_1_metas_118_tag <= cpu_tag_d1;
        end
        if(_zz_637) begin
          ways_1_metas_119_tag <= cpu_tag_d1;
        end
        if(_zz_638) begin
          ways_1_metas_120_tag <= cpu_tag_d1;
        end
        if(_zz_639) begin
          ways_1_metas_121_tag <= cpu_tag_d1;
        end
        if(_zz_640) begin
          ways_1_metas_122_tag <= cpu_tag_d1;
        end
        if(_zz_641) begin
          ways_1_metas_123_tag <= cpu_tag_d1;
        end
        if(_zz_642) begin
          ways_1_metas_124_tag <= cpu_tag_d1;
        end
        if(_zz_643) begin
          ways_1_metas_125_tag <= cpu_tag_d1;
        end
        if(_zz_644) begin
          ways_1_metas_126_tag <= cpu_tag_d1;
        end
        if(_zz_645) begin
          ways_1_metas_127_tag <= cpu_tag_d1;
        end
      end
      if(when_ICache_l230_1) begin
        cpu_cmd_ready_1 <= 1'b0;
      end else begin
        if(when_ICache_l233_1) begin
          cpu_cmd_ready_1 <= 1'b1;
        end
      end
      if(flush_busy) begin
        if(_zz_1034) begin
          ways_2_metas_0_mru <= 1'b0;
        end
        if(_zz_1035) begin
          ways_2_metas_1_mru <= 1'b0;
        end
        if(_zz_1036) begin
          ways_2_metas_2_mru <= 1'b0;
        end
        if(_zz_1037) begin
          ways_2_metas_3_mru <= 1'b0;
        end
        if(_zz_1038) begin
          ways_2_metas_4_mru <= 1'b0;
        end
        if(_zz_1039) begin
          ways_2_metas_5_mru <= 1'b0;
        end
        if(_zz_1040) begin
          ways_2_metas_6_mru <= 1'b0;
        end
        if(_zz_1041) begin
          ways_2_metas_7_mru <= 1'b0;
        end
        if(_zz_1042) begin
          ways_2_metas_8_mru <= 1'b0;
        end
        if(_zz_1043) begin
          ways_2_metas_9_mru <= 1'b0;
        end
        if(_zz_1044) begin
          ways_2_metas_10_mru <= 1'b0;
        end
        if(_zz_1045) begin
          ways_2_metas_11_mru <= 1'b0;
        end
        if(_zz_1046) begin
          ways_2_metas_12_mru <= 1'b0;
        end
        if(_zz_1047) begin
          ways_2_metas_13_mru <= 1'b0;
        end
        if(_zz_1048) begin
          ways_2_metas_14_mru <= 1'b0;
        end
        if(_zz_1049) begin
          ways_2_metas_15_mru <= 1'b0;
        end
        if(_zz_1050) begin
          ways_2_metas_16_mru <= 1'b0;
        end
        if(_zz_1051) begin
          ways_2_metas_17_mru <= 1'b0;
        end
        if(_zz_1052) begin
          ways_2_metas_18_mru <= 1'b0;
        end
        if(_zz_1053) begin
          ways_2_metas_19_mru <= 1'b0;
        end
        if(_zz_1054) begin
          ways_2_metas_20_mru <= 1'b0;
        end
        if(_zz_1055) begin
          ways_2_metas_21_mru <= 1'b0;
        end
        if(_zz_1056) begin
          ways_2_metas_22_mru <= 1'b0;
        end
        if(_zz_1057) begin
          ways_2_metas_23_mru <= 1'b0;
        end
        if(_zz_1058) begin
          ways_2_metas_24_mru <= 1'b0;
        end
        if(_zz_1059) begin
          ways_2_metas_25_mru <= 1'b0;
        end
        if(_zz_1060) begin
          ways_2_metas_26_mru <= 1'b0;
        end
        if(_zz_1061) begin
          ways_2_metas_27_mru <= 1'b0;
        end
        if(_zz_1062) begin
          ways_2_metas_28_mru <= 1'b0;
        end
        if(_zz_1063) begin
          ways_2_metas_29_mru <= 1'b0;
        end
        if(_zz_1064) begin
          ways_2_metas_30_mru <= 1'b0;
        end
        if(_zz_1065) begin
          ways_2_metas_31_mru <= 1'b0;
        end
        if(_zz_1066) begin
          ways_2_metas_32_mru <= 1'b0;
        end
        if(_zz_1067) begin
          ways_2_metas_33_mru <= 1'b0;
        end
        if(_zz_1068) begin
          ways_2_metas_34_mru <= 1'b0;
        end
        if(_zz_1069) begin
          ways_2_metas_35_mru <= 1'b0;
        end
        if(_zz_1070) begin
          ways_2_metas_36_mru <= 1'b0;
        end
        if(_zz_1071) begin
          ways_2_metas_37_mru <= 1'b0;
        end
        if(_zz_1072) begin
          ways_2_metas_38_mru <= 1'b0;
        end
        if(_zz_1073) begin
          ways_2_metas_39_mru <= 1'b0;
        end
        if(_zz_1074) begin
          ways_2_metas_40_mru <= 1'b0;
        end
        if(_zz_1075) begin
          ways_2_metas_41_mru <= 1'b0;
        end
        if(_zz_1076) begin
          ways_2_metas_42_mru <= 1'b0;
        end
        if(_zz_1077) begin
          ways_2_metas_43_mru <= 1'b0;
        end
        if(_zz_1078) begin
          ways_2_metas_44_mru <= 1'b0;
        end
        if(_zz_1079) begin
          ways_2_metas_45_mru <= 1'b0;
        end
        if(_zz_1080) begin
          ways_2_metas_46_mru <= 1'b0;
        end
        if(_zz_1081) begin
          ways_2_metas_47_mru <= 1'b0;
        end
        if(_zz_1082) begin
          ways_2_metas_48_mru <= 1'b0;
        end
        if(_zz_1083) begin
          ways_2_metas_49_mru <= 1'b0;
        end
        if(_zz_1084) begin
          ways_2_metas_50_mru <= 1'b0;
        end
        if(_zz_1085) begin
          ways_2_metas_51_mru <= 1'b0;
        end
        if(_zz_1086) begin
          ways_2_metas_52_mru <= 1'b0;
        end
        if(_zz_1087) begin
          ways_2_metas_53_mru <= 1'b0;
        end
        if(_zz_1088) begin
          ways_2_metas_54_mru <= 1'b0;
        end
        if(_zz_1089) begin
          ways_2_metas_55_mru <= 1'b0;
        end
        if(_zz_1090) begin
          ways_2_metas_56_mru <= 1'b0;
        end
        if(_zz_1091) begin
          ways_2_metas_57_mru <= 1'b0;
        end
        if(_zz_1092) begin
          ways_2_metas_58_mru <= 1'b0;
        end
        if(_zz_1093) begin
          ways_2_metas_59_mru <= 1'b0;
        end
        if(_zz_1094) begin
          ways_2_metas_60_mru <= 1'b0;
        end
        if(_zz_1095) begin
          ways_2_metas_61_mru <= 1'b0;
        end
        if(_zz_1096) begin
          ways_2_metas_62_mru <= 1'b0;
        end
        if(_zz_1097) begin
          ways_2_metas_63_mru <= 1'b0;
        end
        if(_zz_1098) begin
          ways_2_metas_64_mru <= 1'b0;
        end
        if(_zz_1099) begin
          ways_2_metas_65_mru <= 1'b0;
        end
        if(_zz_1100) begin
          ways_2_metas_66_mru <= 1'b0;
        end
        if(_zz_1101) begin
          ways_2_metas_67_mru <= 1'b0;
        end
        if(_zz_1102) begin
          ways_2_metas_68_mru <= 1'b0;
        end
        if(_zz_1103) begin
          ways_2_metas_69_mru <= 1'b0;
        end
        if(_zz_1104) begin
          ways_2_metas_70_mru <= 1'b0;
        end
        if(_zz_1105) begin
          ways_2_metas_71_mru <= 1'b0;
        end
        if(_zz_1106) begin
          ways_2_metas_72_mru <= 1'b0;
        end
        if(_zz_1107) begin
          ways_2_metas_73_mru <= 1'b0;
        end
        if(_zz_1108) begin
          ways_2_metas_74_mru <= 1'b0;
        end
        if(_zz_1109) begin
          ways_2_metas_75_mru <= 1'b0;
        end
        if(_zz_1110) begin
          ways_2_metas_76_mru <= 1'b0;
        end
        if(_zz_1111) begin
          ways_2_metas_77_mru <= 1'b0;
        end
        if(_zz_1112) begin
          ways_2_metas_78_mru <= 1'b0;
        end
        if(_zz_1113) begin
          ways_2_metas_79_mru <= 1'b0;
        end
        if(_zz_1114) begin
          ways_2_metas_80_mru <= 1'b0;
        end
        if(_zz_1115) begin
          ways_2_metas_81_mru <= 1'b0;
        end
        if(_zz_1116) begin
          ways_2_metas_82_mru <= 1'b0;
        end
        if(_zz_1117) begin
          ways_2_metas_83_mru <= 1'b0;
        end
        if(_zz_1118) begin
          ways_2_metas_84_mru <= 1'b0;
        end
        if(_zz_1119) begin
          ways_2_metas_85_mru <= 1'b0;
        end
        if(_zz_1120) begin
          ways_2_metas_86_mru <= 1'b0;
        end
        if(_zz_1121) begin
          ways_2_metas_87_mru <= 1'b0;
        end
        if(_zz_1122) begin
          ways_2_metas_88_mru <= 1'b0;
        end
        if(_zz_1123) begin
          ways_2_metas_89_mru <= 1'b0;
        end
        if(_zz_1124) begin
          ways_2_metas_90_mru <= 1'b0;
        end
        if(_zz_1125) begin
          ways_2_metas_91_mru <= 1'b0;
        end
        if(_zz_1126) begin
          ways_2_metas_92_mru <= 1'b0;
        end
        if(_zz_1127) begin
          ways_2_metas_93_mru <= 1'b0;
        end
        if(_zz_1128) begin
          ways_2_metas_94_mru <= 1'b0;
        end
        if(_zz_1129) begin
          ways_2_metas_95_mru <= 1'b0;
        end
        if(_zz_1130) begin
          ways_2_metas_96_mru <= 1'b0;
        end
        if(_zz_1131) begin
          ways_2_metas_97_mru <= 1'b0;
        end
        if(_zz_1132) begin
          ways_2_metas_98_mru <= 1'b0;
        end
        if(_zz_1133) begin
          ways_2_metas_99_mru <= 1'b0;
        end
        if(_zz_1134) begin
          ways_2_metas_100_mru <= 1'b0;
        end
        if(_zz_1135) begin
          ways_2_metas_101_mru <= 1'b0;
        end
        if(_zz_1136) begin
          ways_2_metas_102_mru <= 1'b0;
        end
        if(_zz_1137) begin
          ways_2_metas_103_mru <= 1'b0;
        end
        if(_zz_1138) begin
          ways_2_metas_104_mru <= 1'b0;
        end
        if(_zz_1139) begin
          ways_2_metas_105_mru <= 1'b0;
        end
        if(_zz_1140) begin
          ways_2_metas_106_mru <= 1'b0;
        end
        if(_zz_1141) begin
          ways_2_metas_107_mru <= 1'b0;
        end
        if(_zz_1142) begin
          ways_2_metas_108_mru <= 1'b0;
        end
        if(_zz_1143) begin
          ways_2_metas_109_mru <= 1'b0;
        end
        if(_zz_1144) begin
          ways_2_metas_110_mru <= 1'b0;
        end
        if(_zz_1145) begin
          ways_2_metas_111_mru <= 1'b0;
        end
        if(_zz_1146) begin
          ways_2_metas_112_mru <= 1'b0;
        end
        if(_zz_1147) begin
          ways_2_metas_113_mru <= 1'b0;
        end
        if(_zz_1148) begin
          ways_2_metas_114_mru <= 1'b0;
        end
        if(_zz_1149) begin
          ways_2_metas_115_mru <= 1'b0;
        end
        if(_zz_1150) begin
          ways_2_metas_116_mru <= 1'b0;
        end
        if(_zz_1151) begin
          ways_2_metas_117_mru <= 1'b0;
        end
        if(_zz_1152) begin
          ways_2_metas_118_mru <= 1'b0;
        end
        if(_zz_1153) begin
          ways_2_metas_119_mru <= 1'b0;
        end
        if(_zz_1154) begin
          ways_2_metas_120_mru <= 1'b0;
        end
        if(_zz_1155) begin
          ways_2_metas_121_mru <= 1'b0;
        end
        if(_zz_1156) begin
          ways_2_metas_122_mru <= 1'b0;
        end
        if(_zz_1157) begin
          ways_2_metas_123_mru <= 1'b0;
        end
        if(_zz_1158) begin
          ways_2_metas_124_mru <= 1'b0;
        end
        if(_zz_1159) begin
          ways_2_metas_125_mru <= 1'b0;
        end
        if(_zz_1160) begin
          ways_2_metas_126_mru <= 1'b0;
        end
        if(_zz_1161) begin
          ways_2_metas_127_mru <= 1'b0;
        end
        if(_zz_1034) begin
          ways_2_metas_0_vld <= 1'b0;
        end
        if(_zz_1035) begin
          ways_2_metas_1_vld <= 1'b0;
        end
        if(_zz_1036) begin
          ways_2_metas_2_vld <= 1'b0;
        end
        if(_zz_1037) begin
          ways_2_metas_3_vld <= 1'b0;
        end
        if(_zz_1038) begin
          ways_2_metas_4_vld <= 1'b0;
        end
        if(_zz_1039) begin
          ways_2_metas_5_vld <= 1'b0;
        end
        if(_zz_1040) begin
          ways_2_metas_6_vld <= 1'b0;
        end
        if(_zz_1041) begin
          ways_2_metas_7_vld <= 1'b0;
        end
        if(_zz_1042) begin
          ways_2_metas_8_vld <= 1'b0;
        end
        if(_zz_1043) begin
          ways_2_metas_9_vld <= 1'b0;
        end
        if(_zz_1044) begin
          ways_2_metas_10_vld <= 1'b0;
        end
        if(_zz_1045) begin
          ways_2_metas_11_vld <= 1'b0;
        end
        if(_zz_1046) begin
          ways_2_metas_12_vld <= 1'b0;
        end
        if(_zz_1047) begin
          ways_2_metas_13_vld <= 1'b0;
        end
        if(_zz_1048) begin
          ways_2_metas_14_vld <= 1'b0;
        end
        if(_zz_1049) begin
          ways_2_metas_15_vld <= 1'b0;
        end
        if(_zz_1050) begin
          ways_2_metas_16_vld <= 1'b0;
        end
        if(_zz_1051) begin
          ways_2_metas_17_vld <= 1'b0;
        end
        if(_zz_1052) begin
          ways_2_metas_18_vld <= 1'b0;
        end
        if(_zz_1053) begin
          ways_2_metas_19_vld <= 1'b0;
        end
        if(_zz_1054) begin
          ways_2_metas_20_vld <= 1'b0;
        end
        if(_zz_1055) begin
          ways_2_metas_21_vld <= 1'b0;
        end
        if(_zz_1056) begin
          ways_2_metas_22_vld <= 1'b0;
        end
        if(_zz_1057) begin
          ways_2_metas_23_vld <= 1'b0;
        end
        if(_zz_1058) begin
          ways_2_metas_24_vld <= 1'b0;
        end
        if(_zz_1059) begin
          ways_2_metas_25_vld <= 1'b0;
        end
        if(_zz_1060) begin
          ways_2_metas_26_vld <= 1'b0;
        end
        if(_zz_1061) begin
          ways_2_metas_27_vld <= 1'b0;
        end
        if(_zz_1062) begin
          ways_2_metas_28_vld <= 1'b0;
        end
        if(_zz_1063) begin
          ways_2_metas_29_vld <= 1'b0;
        end
        if(_zz_1064) begin
          ways_2_metas_30_vld <= 1'b0;
        end
        if(_zz_1065) begin
          ways_2_metas_31_vld <= 1'b0;
        end
        if(_zz_1066) begin
          ways_2_metas_32_vld <= 1'b0;
        end
        if(_zz_1067) begin
          ways_2_metas_33_vld <= 1'b0;
        end
        if(_zz_1068) begin
          ways_2_metas_34_vld <= 1'b0;
        end
        if(_zz_1069) begin
          ways_2_metas_35_vld <= 1'b0;
        end
        if(_zz_1070) begin
          ways_2_metas_36_vld <= 1'b0;
        end
        if(_zz_1071) begin
          ways_2_metas_37_vld <= 1'b0;
        end
        if(_zz_1072) begin
          ways_2_metas_38_vld <= 1'b0;
        end
        if(_zz_1073) begin
          ways_2_metas_39_vld <= 1'b0;
        end
        if(_zz_1074) begin
          ways_2_metas_40_vld <= 1'b0;
        end
        if(_zz_1075) begin
          ways_2_metas_41_vld <= 1'b0;
        end
        if(_zz_1076) begin
          ways_2_metas_42_vld <= 1'b0;
        end
        if(_zz_1077) begin
          ways_2_metas_43_vld <= 1'b0;
        end
        if(_zz_1078) begin
          ways_2_metas_44_vld <= 1'b0;
        end
        if(_zz_1079) begin
          ways_2_metas_45_vld <= 1'b0;
        end
        if(_zz_1080) begin
          ways_2_metas_46_vld <= 1'b0;
        end
        if(_zz_1081) begin
          ways_2_metas_47_vld <= 1'b0;
        end
        if(_zz_1082) begin
          ways_2_metas_48_vld <= 1'b0;
        end
        if(_zz_1083) begin
          ways_2_metas_49_vld <= 1'b0;
        end
        if(_zz_1084) begin
          ways_2_metas_50_vld <= 1'b0;
        end
        if(_zz_1085) begin
          ways_2_metas_51_vld <= 1'b0;
        end
        if(_zz_1086) begin
          ways_2_metas_52_vld <= 1'b0;
        end
        if(_zz_1087) begin
          ways_2_metas_53_vld <= 1'b0;
        end
        if(_zz_1088) begin
          ways_2_metas_54_vld <= 1'b0;
        end
        if(_zz_1089) begin
          ways_2_metas_55_vld <= 1'b0;
        end
        if(_zz_1090) begin
          ways_2_metas_56_vld <= 1'b0;
        end
        if(_zz_1091) begin
          ways_2_metas_57_vld <= 1'b0;
        end
        if(_zz_1092) begin
          ways_2_metas_58_vld <= 1'b0;
        end
        if(_zz_1093) begin
          ways_2_metas_59_vld <= 1'b0;
        end
        if(_zz_1094) begin
          ways_2_metas_60_vld <= 1'b0;
        end
        if(_zz_1095) begin
          ways_2_metas_61_vld <= 1'b0;
        end
        if(_zz_1096) begin
          ways_2_metas_62_vld <= 1'b0;
        end
        if(_zz_1097) begin
          ways_2_metas_63_vld <= 1'b0;
        end
        if(_zz_1098) begin
          ways_2_metas_64_vld <= 1'b0;
        end
        if(_zz_1099) begin
          ways_2_metas_65_vld <= 1'b0;
        end
        if(_zz_1100) begin
          ways_2_metas_66_vld <= 1'b0;
        end
        if(_zz_1101) begin
          ways_2_metas_67_vld <= 1'b0;
        end
        if(_zz_1102) begin
          ways_2_metas_68_vld <= 1'b0;
        end
        if(_zz_1103) begin
          ways_2_metas_69_vld <= 1'b0;
        end
        if(_zz_1104) begin
          ways_2_metas_70_vld <= 1'b0;
        end
        if(_zz_1105) begin
          ways_2_metas_71_vld <= 1'b0;
        end
        if(_zz_1106) begin
          ways_2_metas_72_vld <= 1'b0;
        end
        if(_zz_1107) begin
          ways_2_metas_73_vld <= 1'b0;
        end
        if(_zz_1108) begin
          ways_2_metas_74_vld <= 1'b0;
        end
        if(_zz_1109) begin
          ways_2_metas_75_vld <= 1'b0;
        end
        if(_zz_1110) begin
          ways_2_metas_76_vld <= 1'b0;
        end
        if(_zz_1111) begin
          ways_2_metas_77_vld <= 1'b0;
        end
        if(_zz_1112) begin
          ways_2_metas_78_vld <= 1'b0;
        end
        if(_zz_1113) begin
          ways_2_metas_79_vld <= 1'b0;
        end
        if(_zz_1114) begin
          ways_2_metas_80_vld <= 1'b0;
        end
        if(_zz_1115) begin
          ways_2_metas_81_vld <= 1'b0;
        end
        if(_zz_1116) begin
          ways_2_metas_82_vld <= 1'b0;
        end
        if(_zz_1117) begin
          ways_2_metas_83_vld <= 1'b0;
        end
        if(_zz_1118) begin
          ways_2_metas_84_vld <= 1'b0;
        end
        if(_zz_1119) begin
          ways_2_metas_85_vld <= 1'b0;
        end
        if(_zz_1120) begin
          ways_2_metas_86_vld <= 1'b0;
        end
        if(_zz_1121) begin
          ways_2_metas_87_vld <= 1'b0;
        end
        if(_zz_1122) begin
          ways_2_metas_88_vld <= 1'b0;
        end
        if(_zz_1123) begin
          ways_2_metas_89_vld <= 1'b0;
        end
        if(_zz_1124) begin
          ways_2_metas_90_vld <= 1'b0;
        end
        if(_zz_1125) begin
          ways_2_metas_91_vld <= 1'b0;
        end
        if(_zz_1126) begin
          ways_2_metas_92_vld <= 1'b0;
        end
        if(_zz_1127) begin
          ways_2_metas_93_vld <= 1'b0;
        end
        if(_zz_1128) begin
          ways_2_metas_94_vld <= 1'b0;
        end
        if(_zz_1129) begin
          ways_2_metas_95_vld <= 1'b0;
        end
        if(_zz_1130) begin
          ways_2_metas_96_vld <= 1'b0;
        end
        if(_zz_1131) begin
          ways_2_metas_97_vld <= 1'b0;
        end
        if(_zz_1132) begin
          ways_2_metas_98_vld <= 1'b0;
        end
        if(_zz_1133) begin
          ways_2_metas_99_vld <= 1'b0;
        end
        if(_zz_1134) begin
          ways_2_metas_100_vld <= 1'b0;
        end
        if(_zz_1135) begin
          ways_2_metas_101_vld <= 1'b0;
        end
        if(_zz_1136) begin
          ways_2_metas_102_vld <= 1'b0;
        end
        if(_zz_1137) begin
          ways_2_metas_103_vld <= 1'b0;
        end
        if(_zz_1138) begin
          ways_2_metas_104_vld <= 1'b0;
        end
        if(_zz_1139) begin
          ways_2_metas_105_vld <= 1'b0;
        end
        if(_zz_1140) begin
          ways_2_metas_106_vld <= 1'b0;
        end
        if(_zz_1141) begin
          ways_2_metas_107_vld <= 1'b0;
        end
        if(_zz_1142) begin
          ways_2_metas_108_vld <= 1'b0;
        end
        if(_zz_1143) begin
          ways_2_metas_109_vld <= 1'b0;
        end
        if(_zz_1144) begin
          ways_2_metas_110_vld <= 1'b0;
        end
        if(_zz_1145) begin
          ways_2_metas_111_vld <= 1'b0;
        end
        if(_zz_1146) begin
          ways_2_metas_112_vld <= 1'b0;
        end
        if(_zz_1147) begin
          ways_2_metas_113_vld <= 1'b0;
        end
        if(_zz_1148) begin
          ways_2_metas_114_vld <= 1'b0;
        end
        if(_zz_1149) begin
          ways_2_metas_115_vld <= 1'b0;
        end
        if(_zz_1150) begin
          ways_2_metas_116_vld <= 1'b0;
        end
        if(_zz_1151) begin
          ways_2_metas_117_vld <= 1'b0;
        end
        if(_zz_1152) begin
          ways_2_metas_118_vld <= 1'b0;
        end
        if(_zz_1153) begin
          ways_2_metas_119_vld <= 1'b0;
        end
        if(_zz_1154) begin
          ways_2_metas_120_vld <= 1'b0;
        end
        if(_zz_1155) begin
          ways_2_metas_121_vld <= 1'b0;
        end
        if(_zz_1156) begin
          ways_2_metas_122_vld <= 1'b0;
        end
        if(_zz_1157) begin
          ways_2_metas_123_vld <= 1'b0;
        end
        if(_zz_1158) begin
          ways_2_metas_124_vld <= 1'b0;
        end
        if(_zz_1159) begin
          ways_2_metas_125_vld <= 1'b0;
        end
        if(_zz_1160) begin
          ways_2_metas_126_vld <= 1'b0;
        end
        if(_zz_1161) begin
          ways_2_metas_127_vld <= 1'b0;
        end
      end else begin
        if(when_ICache_l210_2) begin
          if(cache_hit_2) begin
            if(_zz_776) begin
              ways_2_metas_0_mru <= 1'b1;
            end
            if(_zz_777) begin
              ways_2_metas_1_mru <= 1'b1;
            end
            if(_zz_778) begin
              ways_2_metas_2_mru <= 1'b1;
            end
            if(_zz_779) begin
              ways_2_metas_3_mru <= 1'b1;
            end
            if(_zz_780) begin
              ways_2_metas_4_mru <= 1'b1;
            end
            if(_zz_781) begin
              ways_2_metas_5_mru <= 1'b1;
            end
            if(_zz_782) begin
              ways_2_metas_6_mru <= 1'b1;
            end
            if(_zz_783) begin
              ways_2_metas_7_mru <= 1'b1;
            end
            if(_zz_784) begin
              ways_2_metas_8_mru <= 1'b1;
            end
            if(_zz_785) begin
              ways_2_metas_9_mru <= 1'b1;
            end
            if(_zz_786) begin
              ways_2_metas_10_mru <= 1'b1;
            end
            if(_zz_787) begin
              ways_2_metas_11_mru <= 1'b1;
            end
            if(_zz_788) begin
              ways_2_metas_12_mru <= 1'b1;
            end
            if(_zz_789) begin
              ways_2_metas_13_mru <= 1'b1;
            end
            if(_zz_790) begin
              ways_2_metas_14_mru <= 1'b1;
            end
            if(_zz_791) begin
              ways_2_metas_15_mru <= 1'b1;
            end
            if(_zz_792) begin
              ways_2_metas_16_mru <= 1'b1;
            end
            if(_zz_793) begin
              ways_2_metas_17_mru <= 1'b1;
            end
            if(_zz_794) begin
              ways_2_metas_18_mru <= 1'b1;
            end
            if(_zz_795) begin
              ways_2_metas_19_mru <= 1'b1;
            end
            if(_zz_796) begin
              ways_2_metas_20_mru <= 1'b1;
            end
            if(_zz_797) begin
              ways_2_metas_21_mru <= 1'b1;
            end
            if(_zz_798) begin
              ways_2_metas_22_mru <= 1'b1;
            end
            if(_zz_799) begin
              ways_2_metas_23_mru <= 1'b1;
            end
            if(_zz_800) begin
              ways_2_metas_24_mru <= 1'b1;
            end
            if(_zz_801) begin
              ways_2_metas_25_mru <= 1'b1;
            end
            if(_zz_802) begin
              ways_2_metas_26_mru <= 1'b1;
            end
            if(_zz_803) begin
              ways_2_metas_27_mru <= 1'b1;
            end
            if(_zz_804) begin
              ways_2_metas_28_mru <= 1'b1;
            end
            if(_zz_805) begin
              ways_2_metas_29_mru <= 1'b1;
            end
            if(_zz_806) begin
              ways_2_metas_30_mru <= 1'b1;
            end
            if(_zz_807) begin
              ways_2_metas_31_mru <= 1'b1;
            end
            if(_zz_808) begin
              ways_2_metas_32_mru <= 1'b1;
            end
            if(_zz_809) begin
              ways_2_metas_33_mru <= 1'b1;
            end
            if(_zz_810) begin
              ways_2_metas_34_mru <= 1'b1;
            end
            if(_zz_811) begin
              ways_2_metas_35_mru <= 1'b1;
            end
            if(_zz_812) begin
              ways_2_metas_36_mru <= 1'b1;
            end
            if(_zz_813) begin
              ways_2_metas_37_mru <= 1'b1;
            end
            if(_zz_814) begin
              ways_2_metas_38_mru <= 1'b1;
            end
            if(_zz_815) begin
              ways_2_metas_39_mru <= 1'b1;
            end
            if(_zz_816) begin
              ways_2_metas_40_mru <= 1'b1;
            end
            if(_zz_817) begin
              ways_2_metas_41_mru <= 1'b1;
            end
            if(_zz_818) begin
              ways_2_metas_42_mru <= 1'b1;
            end
            if(_zz_819) begin
              ways_2_metas_43_mru <= 1'b1;
            end
            if(_zz_820) begin
              ways_2_metas_44_mru <= 1'b1;
            end
            if(_zz_821) begin
              ways_2_metas_45_mru <= 1'b1;
            end
            if(_zz_822) begin
              ways_2_metas_46_mru <= 1'b1;
            end
            if(_zz_823) begin
              ways_2_metas_47_mru <= 1'b1;
            end
            if(_zz_824) begin
              ways_2_metas_48_mru <= 1'b1;
            end
            if(_zz_825) begin
              ways_2_metas_49_mru <= 1'b1;
            end
            if(_zz_826) begin
              ways_2_metas_50_mru <= 1'b1;
            end
            if(_zz_827) begin
              ways_2_metas_51_mru <= 1'b1;
            end
            if(_zz_828) begin
              ways_2_metas_52_mru <= 1'b1;
            end
            if(_zz_829) begin
              ways_2_metas_53_mru <= 1'b1;
            end
            if(_zz_830) begin
              ways_2_metas_54_mru <= 1'b1;
            end
            if(_zz_831) begin
              ways_2_metas_55_mru <= 1'b1;
            end
            if(_zz_832) begin
              ways_2_metas_56_mru <= 1'b1;
            end
            if(_zz_833) begin
              ways_2_metas_57_mru <= 1'b1;
            end
            if(_zz_834) begin
              ways_2_metas_58_mru <= 1'b1;
            end
            if(_zz_835) begin
              ways_2_metas_59_mru <= 1'b1;
            end
            if(_zz_836) begin
              ways_2_metas_60_mru <= 1'b1;
            end
            if(_zz_837) begin
              ways_2_metas_61_mru <= 1'b1;
            end
            if(_zz_838) begin
              ways_2_metas_62_mru <= 1'b1;
            end
            if(_zz_839) begin
              ways_2_metas_63_mru <= 1'b1;
            end
            if(_zz_840) begin
              ways_2_metas_64_mru <= 1'b1;
            end
            if(_zz_841) begin
              ways_2_metas_65_mru <= 1'b1;
            end
            if(_zz_842) begin
              ways_2_metas_66_mru <= 1'b1;
            end
            if(_zz_843) begin
              ways_2_metas_67_mru <= 1'b1;
            end
            if(_zz_844) begin
              ways_2_metas_68_mru <= 1'b1;
            end
            if(_zz_845) begin
              ways_2_metas_69_mru <= 1'b1;
            end
            if(_zz_846) begin
              ways_2_metas_70_mru <= 1'b1;
            end
            if(_zz_847) begin
              ways_2_metas_71_mru <= 1'b1;
            end
            if(_zz_848) begin
              ways_2_metas_72_mru <= 1'b1;
            end
            if(_zz_849) begin
              ways_2_metas_73_mru <= 1'b1;
            end
            if(_zz_850) begin
              ways_2_metas_74_mru <= 1'b1;
            end
            if(_zz_851) begin
              ways_2_metas_75_mru <= 1'b1;
            end
            if(_zz_852) begin
              ways_2_metas_76_mru <= 1'b1;
            end
            if(_zz_853) begin
              ways_2_metas_77_mru <= 1'b1;
            end
            if(_zz_854) begin
              ways_2_metas_78_mru <= 1'b1;
            end
            if(_zz_855) begin
              ways_2_metas_79_mru <= 1'b1;
            end
            if(_zz_856) begin
              ways_2_metas_80_mru <= 1'b1;
            end
            if(_zz_857) begin
              ways_2_metas_81_mru <= 1'b1;
            end
            if(_zz_858) begin
              ways_2_metas_82_mru <= 1'b1;
            end
            if(_zz_859) begin
              ways_2_metas_83_mru <= 1'b1;
            end
            if(_zz_860) begin
              ways_2_metas_84_mru <= 1'b1;
            end
            if(_zz_861) begin
              ways_2_metas_85_mru <= 1'b1;
            end
            if(_zz_862) begin
              ways_2_metas_86_mru <= 1'b1;
            end
            if(_zz_863) begin
              ways_2_metas_87_mru <= 1'b1;
            end
            if(_zz_864) begin
              ways_2_metas_88_mru <= 1'b1;
            end
            if(_zz_865) begin
              ways_2_metas_89_mru <= 1'b1;
            end
            if(_zz_866) begin
              ways_2_metas_90_mru <= 1'b1;
            end
            if(_zz_867) begin
              ways_2_metas_91_mru <= 1'b1;
            end
            if(_zz_868) begin
              ways_2_metas_92_mru <= 1'b1;
            end
            if(_zz_869) begin
              ways_2_metas_93_mru <= 1'b1;
            end
            if(_zz_870) begin
              ways_2_metas_94_mru <= 1'b1;
            end
            if(_zz_871) begin
              ways_2_metas_95_mru <= 1'b1;
            end
            if(_zz_872) begin
              ways_2_metas_96_mru <= 1'b1;
            end
            if(_zz_873) begin
              ways_2_metas_97_mru <= 1'b1;
            end
            if(_zz_874) begin
              ways_2_metas_98_mru <= 1'b1;
            end
            if(_zz_875) begin
              ways_2_metas_99_mru <= 1'b1;
            end
            if(_zz_876) begin
              ways_2_metas_100_mru <= 1'b1;
            end
            if(_zz_877) begin
              ways_2_metas_101_mru <= 1'b1;
            end
            if(_zz_878) begin
              ways_2_metas_102_mru <= 1'b1;
            end
            if(_zz_879) begin
              ways_2_metas_103_mru <= 1'b1;
            end
            if(_zz_880) begin
              ways_2_metas_104_mru <= 1'b1;
            end
            if(_zz_881) begin
              ways_2_metas_105_mru <= 1'b1;
            end
            if(_zz_882) begin
              ways_2_metas_106_mru <= 1'b1;
            end
            if(_zz_883) begin
              ways_2_metas_107_mru <= 1'b1;
            end
            if(_zz_884) begin
              ways_2_metas_108_mru <= 1'b1;
            end
            if(_zz_885) begin
              ways_2_metas_109_mru <= 1'b1;
            end
            if(_zz_886) begin
              ways_2_metas_110_mru <= 1'b1;
            end
            if(_zz_887) begin
              ways_2_metas_111_mru <= 1'b1;
            end
            if(_zz_888) begin
              ways_2_metas_112_mru <= 1'b1;
            end
            if(_zz_889) begin
              ways_2_metas_113_mru <= 1'b1;
            end
            if(_zz_890) begin
              ways_2_metas_114_mru <= 1'b1;
            end
            if(_zz_891) begin
              ways_2_metas_115_mru <= 1'b1;
            end
            if(_zz_892) begin
              ways_2_metas_116_mru <= 1'b1;
            end
            if(_zz_893) begin
              ways_2_metas_117_mru <= 1'b1;
            end
            if(_zz_894) begin
              ways_2_metas_118_mru <= 1'b1;
            end
            if(_zz_895) begin
              ways_2_metas_119_mru <= 1'b1;
            end
            if(_zz_896) begin
              ways_2_metas_120_mru <= 1'b1;
            end
            if(_zz_897) begin
              ways_2_metas_121_mru <= 1'b1;
            end
            if(_zz_898) begin
              ways_2_metas_122_mru <= 1'b1;
            end
            if(_zz_899) begin
              ways_2_metas_123_mru <= 1'b1;
            end
            if(_zz_900) begin
              ways_2_metas_124_mru <= 1'b1;
            end
            if(_zz_901) begin
              ways_2_metas_125_mru <= 1'b1;
            end
            if(_zz_902) begin
              ways_2_metas_126_mru <= 1'b1;
            end
            if(_zz_903) begin
              ways_2_metas_127_mru <= 1'b1;
            end
          end else begin
            if(_zz_776) begin
              ways_2_metas_0_mru <= 1'b0;
            end
            if(_zz_777) begin
              ways_2_metas_1_mru <= 1'b0;
            end
            if(_zz_778) begin
              ways_2_metas_2_mru <= 1'b0;
            end
            if(_zz_779) begin
              ways_2_metas_3_mru <= 1'b0;
            end
            if(_zz_780) begin
              ways_2_metas_4_mru <= 1'b0;
            end
            if(_zz_781) begin
              ways_2_metas_5_mru <= 1'b0;
            end
            if(_zz_782) begin
              ways_2_metas_6_mru <= 1'b0;
            end
            if(_zz_783) begin
              ways_2_metas_7_mru <= 1'b0;
            end
            if(_zz_784) begin
              ways_2_metas_8_mru <= 1'b0;
            end
            if(_zz_785) begin
              ways_2_metas_9_mru <= 1'b0;
            end
            if(_zz_786) begin
              ways_2_metas_10_mru <= 1'b0;
            end
            if(_zz_787) begin
              ways_2_metas_11_mru <= 1'b0;
            end
            if(_zz_788) begin
              ways_2_metas_12_mru <= 1'b0;
            end
            if(_zz_789) begin
              ways_2_metas_13_mru <= 1'b0;
            end
            if(_zz_790) begin
              ways_2_metas_14_mru <= 1'b0;
            end
            if(_zz_791) begin
              ways_2_metas_15_mru <= 1'b0;
            end
            if(_zz_792) begin
              ways_2_metas_16_mru <= 1'b0;
            end
            if(_zz_793) begin
              ways_2_metas_17_mru <= 1'b0;
            end
            if(_zz_794) begin
              ways_2_metas_18_mru <= 1'b0;
            end
            if(_zz_795) begin
              ways_2_metas_19_mru <= 1'b0;
            end
            if(_zz_796) begin
              ways_2_metas_20_mru <= 1'b0;
            end
            if(_zz_797) begin
              ways_2_metas_21_mru <= 1'b0;
            end
            if(_zz_798) begin
              ways_2_metas_22_mru <= 1'b0;
            end
            if(_zz_799) begin
              ways_2_metas_23_mru <= 1'b0;
            end
            if(_zz_800) begin
              ways_2_metas_24_mru <= 1'b0;
            end
            if(_zz_801) begin
              ways_2_metas_25_mru <= 1'b0;
            end
            if(_zz_802) begin
              ways_2_metas_26_mru <= 1'b0;
            end
            if(_zz_803) begin
              ways_2_metas_27_mru <= 1'b0;
            end
            if(_zz_804) begin
              ways_2_metas_28_mru <= 1'b0;
            end
            if(_zz_805) begin
              ways_2_metas_29_mru <= 1'b0;
            end
            if(_zz_806) begin
              ways_2_metas_30_mru <= 1'b0;
            end
            if(_zz_807) begin
              ways_2_metas_31_mru <= 1'b0;
            end
            if(_zz_808) begin
              ways_2_metas_32_mru <= 1'b0;
            end
            if(_zz_809) begin
              ways_2_metas_33_mru <= 1'b0;
            end
            if(_zz_810) begin
              ways_2_metas_34_mru <= 1'b0;
            end
            if(_zz_811) begin
              ways_2_metas_35_mru <= 1'b0;
            end
            if(_zz_812) begin
              ways_2_metas_36_mru <= 1'b0;
            end
            if(_zz_813) begin
              ways_2_metas_37_mru <= 1'b0;
            end
            if(_zz_814) begin
              ways_2_metas_38_mru <= 1'b0;
            end
            if(_zz_815) begin
              ways_2_metas_39_mru <= 1'b0;
            end
            if(_zz_816) begin
              ways_2_metas_40_mru <= 1'b0;
            end
            if(_zz_817) begin
              ways_2_metas_41_mru <= 1'b0;
            end
            if(_zz_818) begin
              ways_2_metas_42_mru <= 1'b0;
            end
            if(_zz_819) begin
              ways_2_metas_43_mru <= 1'b0;
            end
            if(_zz_820) begin
              ways_2_metas_44_mru <= 1'b0;
            end
            if(_zz_821) begin
              ways_2_metas_45_mru <= 1'b0;
            end
            if(_zz_822) begin
              ways_2_metas_46_mru <= 1'b0;
            end
            if(_zz_823) begin
              ways_2_metas_47_mru <= 1'b0;
            end
            if(_zz_824) begin
              ways_2_metas_48_mru <= 1'b0;
            end
            if(_zz_825) begin
              ways_2_metas_49_mru <= 1'b0;
            end
            if(_zz_826) begin
              ways_2_metas_50_mru <= 1'b0;
            end
            if(_zz_827) begin
              ways_2_metas_51_mru <= 1'b0;
            end
            if(_zz_828) begin
              ways_2_metas_52_mru <= 1'b0;
            end
            if(_zz_829) begin
              ways_2_metas_53_mru <= 1'b0;
            end
            if(_zz_830) begin
              ways_2_metas_54_mru <= 1'b0;
            end
            if(_zz_831) begin
              ways_2_metas_55_mru <= 1'b0;
            end
            if(_zz_832) begin
              ways_2_metas_56_mru <= 1'b0;
            end
            if(_zz_833) begin
              ways_2_metas_57_mru <= 1'b0;
            end
            if(_zz_834) begin
              ways_2_metas_58_mru <= 1'b0;
            end
            if(_zz_835) begin
              ways_2_metas_59_mru <= 1'b0;
            end
            if(_zz_836) begin
              ways_2_metas_60_mru <= 1'b0;
            end
            if(_zz_837) begin
              ways_2_metas_61_mru <= 1'b0;
            end
            if(_zz_838) begin
              ways_2_metas_62_mru <= 1'b0;
            end
            if(_zz_839) begin
              ways_2_metas_63_mru <= 1'b0;
            end
            if(_zz_840) begin
              ways_2_metas_64_mru <= 1'b0;
            end
            if(_zz_841) begin
              ways_2_metas_65_mru <= 1'b0;
            end
            if(_zz_842) begin
              ways_2_metas_66_mru <= 1'b0;
            end
            if(_zz_843) begin
              ways_2_metas_67_mru <= 1'b0;
            end
            if(_zz_844) begin
              ways_2_metas_68_mru <= 1'b0;
            end
            if(_zz_845) begin
              ways_2_metas_69_mru <= 1'b0;
            end
            if(_zz_846) begin
              ways_2_metas_70_mru <= 1'b0;
            end
            if(_zz_847) begin
              ways_2_metas_71_mru <= 1'b0;
            end
            if(_zz_848) begin
              ways_2_metas_72_mru <= 1'b0;
            end
            if(_zz_849) begin
              ways_2_metas_73_mru <= 1'b0;
            end
            if(_zz_850) begin
              ways_2_metas_74_mru <= 1'b0;
            end
            if(_zz_851) begin
              ways_2_metas_75_mru <= 1'b0;
            end
            if(_zz_852) begin
              ways_2_metas_76_mru <= 1'b0;
            end
            if(_zz_853) begin
              ways_2_metas_77_mru <= 1'b0;
            end
            if(_zz_854) begin
              ways_2_metas_78_mru <= 1'b0;
            end
            if(_zz_855) begin
              ways_2_metas_79_mru <= 1'b0;
            end
            if(_zz_856) begin
              ways_2_metas_80_mru <= 1'b0;
            end
            if(_zz_857) begin
              ways_2_metas_81_mru <= 1'b0;
            end
            if(_zz_858) begin
              ways_2_metas_82_mru <= 1'b0;
            end
            if(_zz_859) begin
              ways_2_metas_83_mru <= 1'b0;
            end
            if(_zz_860) begin
              ways_2_metas_84_mru <= 1'b0;
            end
            if(_zz_861) begin
              ways_2_metas_85_mru <= 1'b0;
            end
            if(_zz_862) begin
              ways_2_metas_86_mru <= 1'b0;
            end
            if(_zz_863) begin
              ways_2_metas_87_mru <= 1'b0;
            end
            if(_zz_864) begin
              ways_2_metas_88_mru <= 1'b0;
            end
            if(_zz_865) begin
              ways_2_metas_89_mru <= 1'b0;
            end
            if(_zz_866) begin
              ways_2_metas_90_mru <= 1'b0;
            end
            if(_zz_867) begin
              ways_2_metas_91_mru <= 1'b0;
            end
            if(_zz_868) begin
              ways_2_metas_92_mru <= 1'b0;
            end
            if(_zz_869) begin
              ways_2_metas_93_mru <= 1'b0;
            end
            if(_zz_870) begin
              ways_2_metas_94_mru <= 1'b0;
            end
            if(_zz_871) begin
              ways_2_metas_95_mru <= 1'b0;
            end
            if(_zz_872) begin
              ways_2_metas_96_mru <= 1'b0;
            end
            if(_zz_873) begin
              ways_2_metas_97_mru <= 1'b0;
            end
            if(_zz_874) begin
              ways_2_metas_98_mru <= 1'b0;
            end
            if(_zz_875) begin
              ways_2_metas_99_mru <= 1'b0;
            end
            if(_zz_876) begin
              ways_2_metas_100_mru <= 1'b0;
            end
            if(_zz_877) begin
              ways_2_metas_101_mru <= 1'b0;
            end
            if(_zz_878) begin
              ways_2_metas_102_mru <= 1'b0;
            end
            if(_zz_879) begin
              ways_2_metas_103_mru <= 1'b0;
            end
            if(_zz_880) begin
              ways_2_metas_104_mru <= 1'b0;
            end
            if(_zz_881) begin
              ways_2_metas_105_mru <= 1'b0;
            end
            if(_zz_882) begin
              ways_2_metas_106_mru <= 1'b0;
            end
            if(_zz_883) begin
              ways_2_metas_107_mru <= 1'b0;
            end
            if(_zz_884) begin
              ways_2_metas_108_mru <= 1'b0;
            end
            if(_zz_885) begin
              ways_2_metas_109_mru <= 1'b0;
            end
            if(_zz_886) begin
              ways_2_metas_110_mru <= 1'b0;
            end
            if(_zz_887) begin
              ways_2_metas_111_mru <= 1'b0;
            end
            if(_zz_888) begin
              ways_2_metas_112_mru <= 1'b0;
            end
            if(_zz_889) begin
              ways_2_metas_113_mru <= 1'b0;
            end
            if(_zz_890) begin
              ways_2_metas_114_mru <= 1'b0;
            end
            if(_zz_891) begin
              ways_2_metas_115_mru <= 1'b0;
            end
            if(_zz_892) begin
              ways_2_metas_116_mru <= 1'b0;
            end
            if(_zz_893) begin
              ways_2_metas_117_mru <= 1'b0;
            end
            if(_zz_894) begin
              ways_2_metas_118_mru <= 1'b0;
            end
            if(_zz_895) begin
              ways_2_metas_119_mru <= 1'b0;
            end
            if(_zz_896) begin
              ways_2_metas_120_mru <= 1'b0;
            end
            if(_zz_897) begin
              ways_2_metas_121_mru <= 1'b0;
            end
            if(_zz_898) begin
              ways_2_metas_122_mru <= 1'b0;
            end
            if(_zz_899) begin
              ways_2_metas_123_mru <= 1'b0;
            end
            if(_zz_900) begin
              ways_2_metas_124_mru <= 1'b0;
            end
            if(_zz_901) begin
              ways_2_metas_125_mru <= 1'b0;
            end
            if(_zz_902) begin
              ways_2_metas_126_mru <= 1'b0;
            end
            if(_zz_903) begin
              ways_2_metas_127_mru <= 1'b0;
            end
          end
        end else begin
          if(when_ICache_l217_2) begin
            if(_zz_776) begin
              ways_2_metas_0_mru <= 1'b1;
            end
            if(_zz_777) begin
              ways_2_metas_1_mru <= 1'b1;
            end
            if(_zz_778) begin
              ways_2_metas_2_mru <= 1'b1;
            end
            if(_zz_779) begin
              ways_2_metas_3_mru <= 1'b1;
            end
            if(_zz_780) begin
              ways_2_metas_4_mru <= 1'b1;
            end
            if(_zz_781) begin
              ways_2_metas_5_mru <= 1'b1;
            end
            if(_zz_782) begin
              ways_2_metas_6_mru <= 1'b1;
            end
            if(_zz_783) begin
              ways_2_metas_7_mru <= 1'b1;
            end
            if(_zz_784) begin
              ways_2_metas_8_mru <= 1'b1;
            end
            if(_zz_785) begin
              ways_2_metas_9_mru <= 1'b1;
            end
            if(_zz_786) begin
              ways_2_metas_10_mru <= 1'b1;
            end
            if(_zz_787) begin
              ways_2_metas_11_mru <= 1'b1;
            end
            if(_zz_788) begin
              ways_2_metas_12_mru <= 1'b1;
            end
            if(_zz_789) begin
              ways_2_metas_13_mru <= 1'b1;
            end
            if(_zz_790) begin
              ways_2_metas_14_mru <= 1'b1;
            end
            if(_zz_791) begin
              ways_2_metas_15_mru <= 1'b1;
            end
            if(_zz_792) begin
              ways_2_metas_16_mru <= 1'b1;
            end
            if(_zz_793) begin
              ways_2_metas_17_mru <= 1'b1;
            end
            if(_zz_794) begin
              ways_2_metas_18_mru <= 1'b1;
            end
            if(_zz_795) begin
              ways_2_metas_19_mru <= 1'b1;
            end
            if(_zz_796) begin
              ways_2_metas_20_mru <= 1'b1;
            end
            if(_zz_797) begin
              ways_2_metas_21_mru <= 1'b1;
            end
            if(_zz_798) begin
              ways_2_metas_22_mru <= 1'b1;
            end
            if(_zz_799) begin
              ways_2_metas_23_mru <= 1'b1;
            end
            if(_zz_800) begin
              ways_2_metas_24_mru <= 1'b1;
            end
            if(_zz_801) begin
              ways_2_metas_25_mru <= 1'b1;
            end
            if(_zz_802) begin
              ways_2_metas_26_mru <= 1'b1;
            end
            if(_zz_803) begin
              ways_2_metas_27_mru <= 1'b1;
            end
            if(_zz_804) begin
              ways_2_metas_28_mru <= 1'b1;
            end
            if(_zz_805) begin
              ways_2_metas_29_mru <= 1'b1;
            end
            if(_zz_806) begin
              ways_2_metas_30_mru <= 1'b1;
            end
            if(_zz_807) begin
              ways_2_metas_31_mru <= 1'b1;
            end
            if(_zz_808) begin
              ways_2_metas_32_mru <= 1'b1;
            end
            if(_zz_809) begin
              ways_2_metas_33_mru <= 1'b1;
            end
            if(_zz_810) begin
              ways_2_metas_34_mru <= 1'b1;
            end
            if(_zz_811) begin
              ways_2_metas_35_mru <= 1'b1;
            end
            if(_zz_812) begin
              ways_2_metas_36_mru <= 1'b1;
            end
            if(_zz_813) begin
              ways_2_metas_37_mru <= 1'b1;
            end
            if(_zz_814) begin
              ways_2_metas_38_mru <= 1'b1;
            end
            if(_zz_815) begin
              ways_2_metas_39_mru <= 1'b1;
            end
            if(_zz_816) begin
              ways_2_metas_40_mru <= 1'b1;
            end
            if(_zz_817) begin
              ways_2_metas_41_mru <= 1'b1;
            end
            if(_zz_818) begin
              ways_2_metas_42_mru <= 1'b1;
            end
            if(_zz_819) begin
              ways_2_metas_43_mru <= 1'b1;
            end
            if(_zz_820) begin
              ways_2_metas_44_mru <= 1'b1;
            end
            if(_zz_821) begin
              ways_2_metas_45_mru <= 1'b1;
            end
            if(_zz_822) begin
              ways_2_metas_46_mru <= 1'b1;
            end
            if(_zz_823) begin
              ways_2_metas_47_mru <= 1'b1;
            end
            if(_zz_824) begin
              ways_2_metas_48_mru <= 1'b1;
            end
            if(_zz_825) begin
              ways_2_metas_49_mru <= 1'b1;
            end
            if(_zz_826) begin
              ways_2_metas_50_mru <= 1'b1;
            end
            if(_zz_827) begin
              ways_2_metas_51_mru <= 1'b1;
            end
            if(_zz_828) begin
              ways_2_metas_52_mru <= 1'b1;
            end
            if(_zz_829) begin
              ways_2_metas_53_mru <= 1'b1;
            end
            if(_zz_830) begin
              ways_2_metas_54_mru <= 1'b1;
            end
            if(_zz_831) begin
              ways_2_metas_55_mru <= 1'b1;
            end
            if(_zz_832) begin
              ways_2_metas_56_mru <= 1'b1;
            end
            if(_zz_833) begin
              ways_2_metas_57_mru <= 1'b1;
            end
            if(_zz_834) begin
              ways_2_metas_58_mru <= 1'b1;
            end
            if(_zz_835) begin
              ways_2_metas_59_mru <= 1'b1;
            end
            if(_zz_836) begin
              ways_2_metas_60_mru <= 1'b1;
            end
            if(_zz_837) begin
              ways_2_metas_61_mru <= 1'b1;
            end
            if(_zz_838) begin
              ways_2_metas_62_mru <= 1'b1;
            end
            if(_zz_839) begin
              ways_2_metas_63_mru <= 1'b1;
            end
            if(_zz_840) begin
              ways_2_metas_64_mru <= 1'b1;
            end
            if(_zz_841) begin
              ways_2_metas_65_mru <= 1'b1;
            end
            if(_zz_842) begin
              ways_2_metas_66_mru <= 1'b1;
            end
            if(_zz_843) begin
              ways_2_metas_67_mru <= 1'b1;
            end
            if(_zz_844) begin
              ways_2_metas_68_mru <= 1'b1;
            end
            if(_zz_845) begin
              ways_2_metas_69_mru <= 1'b1;
            end
            if(_zz_846) begin
              ways_2_metas_70_mru <= 1'b1;
            end
            if(_zz_847) begin
              ways_2_metas_71_mru <= 1'b1;
            end
            if(_zz_848) begin
              ways_2_metas_72_mru <= 1'b1;
            end
            if(_zz_849) begin
              ways_2_metas_73_mru <= 1'b1;
            end
            if(_zz_850) begin
              ways_2_metas_74_mru <= 1'b1;
            end
            if(_zz_851) begin
              ways_2_metas_75_mru <= 1'b1;
            end
            if(_zz_852) begin
              ways_2_metas_76_mru <= 1'b1;
            end
            if(_zz_853) begin
              ways_2_metas_77_mru <= 1'b1;
            end
            if(_zz_854) begin
              ways_2_metas_78_mru <= 1'b1;
            end
            if(_zz_855) begin
              ways_2_metas_79_mru <= 1'b1;
            end
            if(_zz_856) begin
              ways_2_metas_80_mru <= 1'b1;
            end
            if(_zz_857) begin
              ways_2_metas_81_mru <= 1'b1;
            end
            if(_zz_858) begin
              ways_2_metas_82_mru <= 1'b1;
            end
            if(_zz_859) begin
              ways_2_metas_83_mru <= 1'b1;
            end
            if(_zz_860) begin
              ways_2_metas_84_mru <= 1'b1;
            end
            if(_zz_861) begin
              ways_2_metas_85_mru <= 1'b1;
            end
            if(_zz_862) begin
              ways_2_metas_86_mru <= 1'b1;
            end
            if(_zz_863) begin
              ways_2_metas_87_mru <= 1'b1;
            end
            if(_zz_864) begin
              ways_2_metas_88_mru <= 1'b1;
            end
            if(_zz_865) begin
              ways_2_metas_89_mru <= 1'b1;
            end
            if(_zz_866) begin
              ways_2_metas_90_mru <= 1'b1;
            end
            if(_zz_867) begin
              ways_2_metas_91_mru <= 1'b1;
            end
            if(_zz_868) begin
              ways_2_metas_92_mru <= 1'b1;
            end
            if(_zz_869) begin
              ways_2_metas_93_mru <= 1'b1;
            end
            if(_zz_870) begin
              ways_2_metas_94_mru <= 1'b1;
            end
            if(_zz_871) begin
              ways_2_metas_95_mru <= 1'b1;
            end
            if(_zz_872) begin
              ways_2_metas_96_mru <= 1'b1;
            end
            if(_zz_873) begin
              ways_2_metas_97_mru <= 1'b1;
            end
            if(_zz_874) begin
              ways_2_metas_98_mru <= 1'b1;
            end
            if(_zz_875) begin
              ways_2_metas_99_mru <= 1'b1;
            end
            if(_zz_876) begin
              ways_2_metas_100_mru <= 1'b1;
            end
            if(_zz_877) begin
              ways_2_metas_101_mru <= 1'b1;
            end
            if(_zz_878) begin
              ways_2_metas_102_mru <= 1'b1;
            end
            if(_zz_879) begin
              ways_2_metas_103_mru <= 1'b1;
            end
            if(_zz_880) begin
              ways_2_metas_104_mru <= 1'b1;
            end
            if(_zz_881) begin
              ways_2_metas_105_mru <= 1'b1;
            end
            if(_zz_882) begin
              ways_2_metas_106_mru <= 1'b1;
            end
            if(_zz_883) begin
              ways_2_metas_107_mru <= 1'b1;
            end
            if(_zz_884) begin
              ways_2_metas_108_mru <= 1'b1;
            end
            if(_zz_885) begin
              ways_2_metas_109_mru <= 1'b1;
            end
            if(_zz_886) begin
              ways_2_metas_110_mru <= 1'b1;
            end
            if(_zz_887) begin
              ways_2_metas_111_mru <= 1'b1;
            end
            if(_zz_888) begin
              ways_2_metas_112_mru <= 1'b1;
            end
            if(_zz_889) begin
              ways_2_metas_113_mru <= 1'b1;
            end
            if(_zz_890) begin
              ways_2_metas_114_mru <= 1'b1;
            end
            if(_zz_891) begin
              ways_2_metas_115_mru <= 1'b1;
            end
            if(_zz_892) begin
              ways_2_metas_116_mru <= 1'b1;
            end
            if(_zz_893) begin
              ways_2_metas_117_mru <= 1'b1;
            end
            if(_zz_894) begin
              ways_2_metas_118_mru <= 1'b1;
            end
            if(_zz_895) begin
              ways_2_metas_119_mru <= 1'b1;
            end
            if(_zz_896) begin
              ways_2_metas_120_mru <= 1'b1;
            end
            if(_zz_897) begin
              ways_2_metas_121_mru <= 1'b1;
            end
            if(_zz_898) begin
              ways_2_metas_122_mru <= 1'b1;
            end
            if(_zz_899) begin
              ways_2_metas_123_mru <= 1'b1;
            end
            if(_zz_900) begin
              ways_2_metas_124_mru <= 1'b1;
            end
            if(_zz_901) begin
              ways_2_metas_125_mru <= 1'b1;
            end
            if(_zz_902) begin
              ways_2_metas_126_mru <= 1'b1;
            end
            if(_zz_903) begin
              ways_2_metas_127_mru <= 1'b1;
            end
          end else begin
            if(when_ICache_l220_2) begin
              if(_zz_905) begin
                ways_2_metas_0_vld <= 1'b1;
              end
              if(_zz_906) begin
                ways_2_metas_1_vld <= 1'b1;
              end
              if(_zz_907) begin
                ways_2_metas_2_vld <= 1'b1;
              end
              if(_zz_908) begin
                ways_2_metas_3_vld <= 1'b1;
              end
              if(_zz_909) begin
                ways_2_metas_4_vld <= 1'b1;
              end
              if(_zz_910) begin
                ways_2_metas_5_vld <= 1'b1;
              end
              if(_zz_911) begin
                ways_2_metas_6_vld <= 1'b1;
              end
              if(_zz_912) begin
                ways_2_metas_7_vld <= 1'b1;
              end
              if(_zz_913) begin
                ways_2_metas_8_vld <= 1'b1;
              end
              if(_zz_914) begin
                ways_2_metas_9_vld <= 1'b1;
              end
              if(_zz_915) begin
                ways_2_metas_10_vld <= 1'b1;
              end
              if(_zz_916) begin
                ways_2_metas_11_vld <= 1'b1;
              end
              if(_zz_917) begin
                ways_2_metas_12_vld <= 1'b1;
              end
              if(_zz_918) begin
                ways_2_metas_13_vld <= 1'b1;
              end
              if(_zz_919) begin
                ways_2_metas_14_vld <= 1'b1;
              end
              if(_zz_920) begin
                ways_2_metas_15_vld <= 1'b1;
              end
              if(_zz_921) begin
                ways_2_metas_16_vld <= 1'b1;
              end
              if(_zz_922) begin
                ways_2_metas_17_vld <= 1'b1;
              end
              if(_zz_923) begin
                ways_2_metas_18_vld <= 1'b1;
              end
              if(_zz_924) begin
                ways_2_metas_19_vld <= 1'b1;
              end
              if(_zz_925) begin
                ways_2_metas_20_vld <= 1'b1;
              end
              if(_zz_926) begin
                ways_2_metas_21_vld <= 1'b1;
              end
              if(_zz_927) begin
                ways_2_metas_22_vld <= 1'b1;
              end
              if(_zz_928) begin
                ways_2_metas_23_vld <= 1'b1;
              end
              if(_zz_929) begin
                ways_2_metas_24_vld <= 1'b1;
              end
              if(_zz_930) begin
                ways_2_metas_25_vld <= 1'b1;
              end
              if(_zz_931) begin
                ways_2_metas_26_vld <= 1'b1;
              end
              if(_zz_932) begin
                ways_2_metas_27_vld <= 1'b1;
              end
              if(_zz_933) begin
                ways_2_metas_28_vld <= 1'b1;
              end
              if(_zz_934) begin
                ways_2_metas_29_vld <= 1'b1;
              end
              if(_zz_935) begin
                ways_2_metas_30_vld <= 1'b1;
              end
              if(_zz_936) begin
                ways_2_metas_31_vld <= 1'b1;
              end
              if(_zz_937) begin
                ways_2_metas_32_vld <= 1'b1;
              end
              if(_zz_938) begin
                ways_2_metas_33_vld <= 1'b1;
              end
              if(_zz_939) begin
                ways_2_metas_34_vld <= 1'b1;
              end
              if(_zz_940) begin
                ways_2_metas_35_vld <= 1'b1;
              end
              if(_zz_941) begin
                ways_2_metas_36_vld <= 1'b1;
              end
              if(_zz_942) begin
                ways_2_metas_37_vld <= 1'b1;
              end
              if(_zz_943) begin
                ways_2_metas_38_vld <= 1'b1;
              end
              if(_zz_944) begin
                ways_2_metas_39_vld <= 1'b1;
              end
              if(_zz_945) begin
                ways_2_metas_40_vld <= 1'b1;
              end
              if(_zz_946) begin
                ways_2_metas_41_vld <= 1'b1;
              end
              if(_zz_947) begin
                ways_2_metas_42_vld <= 1'b1;
              end
              if(_zz_948) begin
                ways_2_metas_43_vld <= 1'b1;
              end
              if(_zz_949) begin
                ways_2_metas_44_vld <= 1'b1;
              end
              if(_zz_950) begin
                ways_2_metas_45_vld <= 1'b1;
              end
              if(_zz_951) begin
                ways_2_metas_46_vld <= 1'b1;
              end
              if(_zz_952) begin
                ways_2_metas_47_vld <= 1'b1;
              end
              if(_zz_953) begin
                ways_2_metas_48_vld <= 1'b1;
              end
              if(_zz_954) begin
                ways_2_metas_49_vld <= 1'b1;
              end
              if(_zz_955) begin
                ways_2_metas_50_vld <= 1'b1;
              end
              if(_zz_956) begin
                ways_2_metas_51_vld <= 1'b1;
              end
              if(_zz_957) begin
                ways_2_metas_52_vld <= 1'b1;
              end
              if(_zz_958) begin
                ways_2_metas_53_vld <= 1'b1;
              end
              if(_zz_959) begin
                ways_2_metas_54_vld <= 1'b1;
              end
              if(_zz_960) begin
                ways_2_metas_55_vld <= 1'b1;
              end
              if(_zz_961) begin
                ways_2_metas_56_vld <= 1'b1;
              end
              if(_zz_962) begin
                ways_2_metas_57_vld <= 1'b1;
              end
              if(_zz_963) begin
                ways_2_metas_58_vld <= 1'b1;
              end
              if(_zz_964) begin
                ways_2_metas_59_vld <= 1'b1;
              end
              if(_zz_965) begin
                ways_2_metas_60_vld <= 1'b1;
              end
              if(_zz_966) begin
                ways_2_metas_61_vld <= 1'b1;
              end
              if(_zz_967) begin
                ways_2_metas_62_vld <= 1'b1;
              end
              if(_zz_968) begin
                ways_2_metas_63_vld <= 1'b1;
              end
              if(_zz_969) begin
                ways_2_metas_64_vld <= 1'b1;
              end
              if(_zz_970) begin
                ways_2_metas_65_vld <= 1'b1;
              end
              if(_zz_971) begin
                ways_2_metas_66_vld <= 1'b1;
              end
              if(_zz_972) begin
                ways_2_metas_67_vld <= 1'b1;
              end
              if(_zz_973) begin
                ways_2_metas_68_vld <= 1'b1;
              end
              if(_zz_974) begin
                ways_2_metas_69_vld <= 1'b1;
              end
              if(_zz_975) begin
                ways_2_metas_70_vld <= 1'b1;
              end
              if(_zz_976) begin
                ways_2_metas_71_vld <= 1'b1;
              end
              if(_zz_977) begin
                ways_2_metas_72_vld <= 1'b1;
              end
              if(_zz_978) begin
                ways_2_metas_73_vld <= 1'b1;
              end
              if(_zz_979) begin
                ways_2_metas_74_vld <= 1'b1;
              end
              if(_zz_980) begin
                ways_2_metas_75_vld <= 1'b1;
              end
              if(_zz_981) begin
                ways_2_metas_76_vld <= 1'b1;
              end
              if(_zz_982) begin
                ways_2_metas_77_vld <= 1'b1;
              end
              if(_zz_983) begin
                ways_2_metas_78_vld <= 1'b1;
              end
              if(_zz_984) begin
                ways_2_metas_79_vld <= 1'b1;
              end
              if(_zz_985) begin
                ways_2_metas_80_vld <= 1'b1;
              end
              if(_zz_986) begin
                ways_2_metas_81_vld <= 1'b1;
              end
              if(_zz_987) begin
                ways_2_metas_82_vld <= 1'b1;
              end
              if(_zz_988) begin
                ways_2_metas_83_vld <= 1'b1;
              end
              if(_zz_989) begin
                ways_2_metas_84_vld <= 1'b1;
              end
              if(_zz_990) begin
                ways_2_metas_85_vld <= 1'b1;
              end
              if(_zz_991) begin
                ways_2_metas_86_vld <= 1'b1;
              end
              if(_zz_992) begin
                ways_2_metas_87_vld <= 1'b1;
              end
              if(_zz_993) begin
                ways_2_metas_88_vld <= 1'b1;
              end
              if(_zz_994) begin
                ways_2_metas_89_vld <= 1'b1;
              end
              if(_zz_995) begin
                ways_2_metas_90_vld <= 1'b1;
              end
              if(_zz_996) begin
                ways_2_metas_91_vld <= 1'b1;
              end
              if(_zz_997) begin
                ways_2_metas_92_vld <= 1'b1;
              end
              if(_zz_998) begin
                ways_2_metas_93_vld <= 1'b1;
              end
              if(_zz_999) begin
                ways_2_metas_94_vld <= 1'b1;
              end
              if(_zz_1000) begin
                ways_2_metas_95_vld <= 1'b1;
              end
              if(_zz_1001) begin
                ways_2_metas_96_vld <= 1'b1;
              end
              if(_zz_1002) begin
                ways_2_metas_97_vld <= 1'b1;
              end
              if(_zz_1003) begin
                ways_2_metas_98_vld <= 1'b1;
              end
              if(_zz_1004) begin
                ways_2_metas_99_vld <= 1'b1;
              end
              if(_zz_1005) begin
                ways_2_metas_100_vld <= 1'b1;
              end
              if(_zz_1006) begin
                ways_2_metas_101_vld <= 1'b1;
              end
              if(_zz_1007) begin
                ways_2_metas_102_vld <= 1'b1;
              end
              if(_zz_1008) begin
                ways_2_metas_103_vld <= 1'b1;
              end
              if(_zz_1009) begin
                ways_2_metas_104_vld <= 1'b1;
              end
              if(_zz_1010) begin
                ways_2_metas_105_vld <= 1'b1;
              end
              if(_zz_1011) begin
                ways_2_metas_106_vld <= 1'b1;
              end
              if(_zz_1012) begin
                ways_2_metas_107_vld <= 1'b1;
              end
              if(_zz_1013) begin
                ways_2_metas_108_vld <= 1'b1;
              end
              if(_zz_1014) begin
                ways_2_metas_109_vld <= 1'b1;
              end
              if(_zz_1015) begin
                ways_2_metas_110_vld <= 1'b1;
              end
              if(_zz_1016) begin
                ways_2_metas_111_vld <= 1'b1;
              end
              if(_zz_1017) begin
                ways_2_metas_112_vld <= 1'b1;
              end
              if(_zz_1018) begin
                ways_2_metas_113_vld <= 1'b1;
              end
              if(_zz_1019) begin
                ways_2_metas_114_vld <= 1'b1;
              end
              if(_zz_1020) begin
                ways_2_metas_115_vld <= 1'b1;
              end
              if(_zz_1021) begin
                ways_2_metas_116_vld <= 1'b1;
              end
              if(_zz_1022) begin
                ways_2_metas_117_vld <= 1'b1;
              end
              if(_zz_1023) begin
                ways_2_metas_118_vld <= 1'b1;
              end
              if(_zz_1024) begin
                ways_2_metas_119_vld <= 1'b1;
              end
              if(_zz_1025) begin
                ways_2_metas_120_vld <= 1'b1;
              end
              if(_zz_1026) begin
                ways_2_metas_121_vld <= 1'b1;
              end
              if(_zz_1027) begin
                ways_2_metas_122_vld <= 1'b1;
              end
              if(_zz_1028) begin
                ways_2_metas_123_vld <= 1'b1;
              end
              if(_zz_1029) begin
                ways_2_metas_124_vld <= 1'b1;
              end
              if(_zz_1030) begin
                ways_2_metas_125_vld <= 1'b1;
              end
              if(_zz_1031) begin
                ways_2_metas_126_vld <= 1'b1;
              end
              if(_zz_1032) begin
                ways_2_metas_127_vld <= 1'b1;
              end
            end
          end
        end
      end
      if(when_ICache_l225_2) begin
        if(_zz_905) begin
          ways_2_metas_0_tag <= cpu_tag_d1;
        end
        if(_zz_906) begin
          ways_2_metas_1_tag <= cpu_tag_d1;
        end
        if(_zz_907) begin
          ways_2_metas_2_tag <= cpu_tag_d1;
        end
        if(_zz_908) begin
          ways_2_metas_3_tag <= cpu_tag_d1;
        end
        if(_zz_909) begin
          ways_2_metas_4_tag <= cpu_tag_d1;
        end
        if(_zz_910) begin
          ways_2_metas_5_tag <= cpu_tag_d1;
        end
        if(_zz_911) begin
          ways_2_metas_6_tag <= cpu_tag_d1;
        end
        if(_zz_912) begin
          ways_2_metas_7_tag <= cpu_tag_d1;
        end
        if(_zz_913) begin
          ways_2_metas_8_tag <= cpu_tag_d1;
        end
        if(_zz_914) begin
          ways_2_metas_9_tag <= cpu_tag_d1;
        end
        if(_zz_915) begin
          ways_2_metas_10_tag <= cpu_tag_d1;
        end
        if(_zz_916) begin
          ways_2_metas_11_tag <= cpu_tag_d1;
        end
        if(_zz_917) begin
          ways_2_metas_12_tag <= cpu_tag_d1;
        end
        if(_zz_918) begin
          ways_2_metas_13_tag <= cpu_tag_d1;
        end
        if(_zz_919) begin
          ways_2_metas_14_tag <= cpu_tag_d1;
        end
        if(_zz_920) begin
          ways_2_metas_15_tag <= cpu_tag_d1;
        end
        if(_zz_921) begin
          ways_2_metas_16_tag <= cpu_tag_d1;
        end
        if(_zz_922) begin
          ways_2_metas_17_tag <= cpu_tag_d1;
        end
        if(_zz_923) begin
          ways_2_metas_18_tag <= cpu_tag_d1;
        end
        if(_zz_924) begin
          ways_2_metas_19_tag <= cpu_tag_d1;
        end
        if(_zz_925) begin
          ways_2_metas_20_tag <= cpu_tag_d1;
        end
        if(_zz_926) begin
          ways_2_metas_21_tag <= cpu_tag_d1;
        end
        if(_zz_927) begin
          ways_2_metas_22_tag <= cpu_tag_d1;
        end
        if(_zz_928) begin
          ways_2_metas_23_tag <= cpu_tag_d1;
        end
        if(_zz_929) begin
          ways_2_metas_24_tag <= cpu_tag_d1;
        end
        if(_zz_930) begin
          ways_2_metas_25_tag <= cpu_tag_d1;
        end
        if(_zz_931) begin
          ways_2_metas_26_tag <= cpu_tag_d1;
        end
        if(_zz_932) begin
          ways_2_metas_27_tag <= cpu_tag_d1;
        end
        if(_zz_933) begin
          ways_2_metas_28_tag <= cpu_tag_d1;
        end
        if(_zz_934) begin
          ways_2_metas_29_tag <= cpu_tag_d1;
        end
        if(_zz_935) begin
          ways_2_metas_30_tag <= cpu_tag_d1;
        end
        if(_zz_936) begin
          ways_2_metas_31_tag <= cpu_tag_d1;
        end
        if(_zz_937) begin
          ways_2_metas_32_tag <= cpu_tag_d1;
        end
        if(_zz_938) begin
          ways_2_metas_33_tag <= cpu_tag_d1;
        end
        if(_zz_939) begin
          ways_2_metas_34_tag <= cpu_tag_d1;
        end
        if(_zz_940) begin
          ways_2_metas_35_tag <= cpu_tag_d1;
        end
        if(_zz_941) begin
          ways_2_metas_36_tag <= cpu_tag_d1;
        end
        if(_zz_942) begin
          ways_2_metas_37_tag <= cpu_tag_d1;
        end
        if(_zz_943) begin
          ways_2_metas_38_tag <= cpu_tag_d1;
        end
        if(_zz_944) begin
          ways_2_metas_39_tag <= cpu_tag_d1;
        end
        if(_zz_945) begin
          ways_2_metas_40_tag <= cpu_tag_d1;
        end
        if(_zz_946) begin
          ways_2_metas_41_tag <= cpu_tag_d1;
        end
        if(_zz_947) begin
          ways_2_metas_42_tag <= cpu_tag_d1;
        end
        if(_zz_948) begin
          ways_2_metas_43_tag <= cpu_tag_d1;
        end
        if(_zz_949) begin
          ways_2_metas_44_tag <= cpu_tag_d1;
        end
        if(_zz_950) begin
          ways_2_metas_45_tag <= cpu_tag_d1;
        end
        if(_zz_951) begin
          ways_2_metas_46_tag <= cpu_tag_d1;
        end
        if(_zz_952) begin
          ways_2_metas_47_tag <= cpu_tag_d1;
        end
        if(_zz_953) begin
          ways_2_metas_48_tag <= cpu_tag_d1;
        end
        if(_zz_954) begin
          ways_2_metas_49_tag <= cpu_tag_d1;
        end
        if(_zz_955) begin
          ways_2_metas_50_tag <= cpu_tag_d1;
        end
        if(_zz_956) begin
          ways_2_metas_51_tag <= cpu_tag_d1;
        end
        if(_zz_957) begin
          ways_2_metas_52_tag <= cpu_tag_d1;
        end
        if(_zz_958) begin
          ways_2_metas_53_tag <= cpu_tag_d1;
        end
        if(_zz_959) begin
          ways_2_metas_54_tag <= cpu_tag_d1;
        end
        if(_zz_960) begin
          ways_2_metas_55_tag <= cpu_tag_d1;
        end
        if(_zz_961) begin
          ways_2_metas_56_tag <= cpu_tag_d1;
        end
        if(_zz_962) begin
          ways_2_metas_57_tag <= cpu_tag_d1;
        end
        if(_zz_963) begin
          ways_2_metas_58_tag <= cpu_tag_d1;
        end
        if(_zz_964) begin
          ways_2_metas_59_tag <= cpu_tag_d1;
        end
        if(_zz_965) begin
          ways_2_metas_60_tag <= cpu_tag_d1;
        end
        if(_zz_966) begin
          ways_2_metas_61_tag <= cpu_tag_d1;
        end
        if(_zz_967) begin
          ways_2_metas_62_tag <= cpu_tag_d1;
        end
        if(_zz_968) begin
          ways_2_metas_63_tag <= cpu_tag_d1;
        end
        if(_zz_969) begin
          ways_2_metas_64_tag <= cpu_tag_d1;
        end
        if(_zz_970) begin
          ways_2_metas_65_tag <= cpu_tag_d1;
        end
        if(_zz_971) begin
          ways_2_metas_66_tag <= cpu_tag_d1;
        end
        if(_zz_972) begin
          ways_2_metas_67_tag <= cpu_tag_d1;
        end
        if(_zz_973) begin
          ways_2_metas_68_tag <= cpu_tag_d1;
        end
        if(_zz_974) begin
          ways_2_metas_69_tag <= cpu_tag_d1;
        end
        if(_zz_975) begin
          ways_2_metas_70_tag <= cpu_tag_d1;
        end
        if(_zz_976) begin
          ways_2_metas_71_tag <= cpu_tag_d1;
        end
        if(_zz_977) begin
          ways_2_metas_72_tag <= cpu_tag_d1;
        end
        if(_zz_978) begin
          ways_2_metas_73_tag <= cpu_tag_d1;
        end
        if(_zz_979) begin
          ways_2_metas_74_tag <= cpu_tag_d1;
        end
        if(_zz_980) begin
          ways_2_metas_75_tag <= cpu_tag_d1;
        end
        if(_zz_981) begin
          ways_2_metas_76_tag <= cpu_tag_d1;
        end
        if(_zz_982) begin
          ways_2_metas_77_tag <= cpu_tag_d1;
        end
        if(_zz_983) begin
          ways_2_metas_78_tag <= cpu_tag_d1;
        end
        if(_zz_984) begin
          ways_2_metas_79_tag <= cpu_tag_d1;
        end
        if(_zz_985) begin
          ways_2_metas_80_tag <= cpu_tag_d1;
        end
        if(_zz_986) begin
          ways_2_metas_81_tag <= cpu_tag_d1;
        end
        if(_zz_987) begin
          ways_2_metas_82_tag <= cpu_tag_d1;
        end
        if(_zz_988) begin
          ways_2_metas_83_tag <= cpu_tag_d1;
        end
        if(_zz_989) begin
          ways_2_metas_84_tag <= cpu_tag_d1;
        end
        if(_zz_990) begin
          ways_2_metas_85_tag <= cpu_tag_d1;
        end
        if(_zz_991) begin
          ways_2_metas_86_tag <= cpu_tag_d1;
        end
        if(_zz_992) begin
          ways_2_metas_87_tag <= cpu_tag_d1;
        end
        if(_zz_993) begin
          ways_2_metas_88_tag <= cpu_tag_d1;
        end
        if(_zz_994) begin
          ways_2_metas_89_tag <= cpu_tag_d1;
        end
        if(_zz_995) begin
          ways_2_metas_90_tag <= cpu_tag_d1;
        end
        if(_zz_996) begin
          ways_2_metas_91_tag <= cpu_tag_d1;
        end
        if(_zz_997) begin
          ways_2_metas_92_tag <= cpu_tag_d1;
        end
        if(_zz_998) begin
          ways_2_metas_93_tag <= cpu_tag_d1;
        end
        if(_zz_999) begin
          ways_2_metas_94_tag <= cpu_tag_d1;
        end
        if(_zz_1000) begin
          ways_2_metas_95_tag <= cpu_tag_d1;
        end
        if(_zz_1001) begin
          ways_2_metas_96_tag <= cpu_tag_d1;
        end
        if(_zz_1002) begin
          ways_2_metas_97_tag <= cpu_tag_d1;
        end
        if(_zz_1003) begin
          ways_2_metas_98_tag <= cpu_tag_d1;
        end
        if(_zz_1004) begin
          ways_2_metas_99_tag <= cpu_tag_d1;
        end
        if(_zz_1005) begin
          ways_2_metas_100_tag <= cpu_tag_d1;
        end
        if(_zz_1006) begin
          ways_2_metas_101_tag <= cpu_tag_d1;
        end
        if(_zz_1007) begin
          ways_2_metas_102_tag <= cpu_tag_d1;
        end
        if(_zz_1008) begin
          ways_2_metas_103_tag <= cpu_tag_d1;
        end
        if(_zz_1009) begin
          ways_2_metas_104_tag <= cpu_tag_d1;
        end
        if(_zz_1010) begin
          ways_2_metas_105_tag <= cpu_tag_d1;
        end
        if(_zz_1011) begin
          ways_2_metas_106_tag <= cpu_tag_d1;
        end
        if(_zz_1012) begin
          ways_2_metas_107_tag <= cpu_tag_d1;
        end
        if(_zz_1013) begin
          ways_2_metas_108_tag <= cpu_tag_d1;
        end
        if(_zz_1014) begin
          ways_2_metas_109_tag <= cpu_tag_d1;
        end
        if(_zz_1015) begin
          ways_2_metas_110_tag <= cpu_tag_d1;
        end
        if(_zz_1016) begin
          ways_2_metas_111_tag <= cpu_tag_d1;
        end
        if(_zz_1017) begin
          ways_2_metas_112_tag <= cpu_tag_d1;
        end
        if(_zz_1018) begin
          ways_2_metas_113_tag <= cpu_tag_d1;
        end
        if(_zz_1019) begin
          ways_2_metas_114_tag <= cpu_tag_d1;
        end
        if(_zz_1020) begin
          ways_2_metas_115_tag <= cpu_tag_d1;
        end
        if(_zz_1021) begin
          ways_2_metas_116_tag <= cpu_tag_d1;
        end
        if(_zz_1022) begin
          ways_2_metas_117_tag <= cpu_tag_d1;
        end
        if(_zz_1023) begin
          ways_2_metas_118_tag <= cpu_tag_d1;
        end
        if(_zz_1024) begin
          ways_2_metas_119_tag <= cpu_tag_d1;
        end
        if(_zz_1025) begin
          ways_2_metas_120_tag <= cpu_tag_d1;
        end
        if(_zz_1026) begin
          ways_2_metas_121_tag <= cpu_tag_d1;
        end
        if(_zz_1027) begin
          ways_2_metas_122_tag <= cpu_tag_d1;
        end
        if(_zz_1028) begin
          ways_2_metas_123_tag <= cpu_tag_d1;
        end
        if(_zz_1029) begin
          ways_2_metas_124_tag <= cpu_tag_d1;
        end
        if(_zz_1030) begin
          ways_2_metas_125_tag <= cpu_tag_d1;
        end
        if(_zz_1031) begin
          ways_2_metas_126_tag <= cpu_tag_d1;
        end
        if(_zz_1032) begin
          ways_2_metas_127_tag <= cpu_tag_d1;
        end
      end
      if(when_ICache_l230_2) begin
        cpu_cmd_ready_1 <= 1'b0;
      end else begin
        if(when_ICache_l233_2) begin
          cpu_cmd_ready_1 <= 1'b1;
        end
      end
      if(flush_busy) begin
        if(_zz_1421) begin
          ways_3_metas_0_mru <= 1'b0;
        end
        if(_zz_1422) begin
          ways_3_metas_1_mru <= 1'b0;
        end
        if(_zz_1423) begin
          ways_3_metas_2_mru <= 1'b0;
        end
        if(_zz_1424) begin
          ways_3_metas_3_mru <= 1'b0;
        end
        if(_zz_1425) begin
          ways_3_metas_4_mru <= 1'b0;
        end
        if(_zz_1426) begin
          ways_3_metas_5_mru <= 1'b0;
        end
        if(_zz_1427) begin
          ways_3_metas_6_mru <= 1'b0;
        end
        if(_zz_1428) begin
          ways_3_metas_7_mru <= 1'b0;
        end
        if(_zz_1429) begin
          ways_3_metas_8_mru <= 1'b0;
        end
        if(_zz_1430) begin
          ways_3_metas_9_mru <= 1'b0;
        end
        if(_zz_1431) begin
          ways_3_metas_10_mru <= 1'b0;
        end
        if(_zz_1432) begin
          ways_3_metas_11_mru <= 1'b0;
        end
        if(_zz_1433) begin
          ways_3_metas_12_mru <= 1'b0;
        end
        if(_zz_1434) begin
          ways_3_metas_13_mru <= 1'b0;
        end
        if(_zz_1435) begin
          ways_3_metas_14_mru <= 1'b0;
        end
        if(_zz_1436) begin
          ways_3_metas_15_mru <= 1'b0;
        end
        if(_zz_1437) begin
          ways_3_metas_16_mru <= 1'b0;
        end
        if(_zz_1438) begin
          ways_3_metas_17_mru <= 1'b0;
        end
        if(_zz_1439) begin
          ways_3_metas_18_mru <= 1'b0;
        end
        if(_zz_1440) begin
          ways_3_metas_19_mru <= 1'b0;
        end
        if(_zz_1441) begin
          ways_3_metas_20_mru <= 1'b0;
        end
        if(_zz_1442) begin
          ways_3_metas_21_mru <= 1'b0;
        end
        if(_zz_1443) begin
          ways_3_metas_22_mru <= 1'b0;
        end
        if(_zz_1444) begin
          ways_3_metas_23_mru <= 1'b0;
        end
        if(_zz_1445) begin
          ways_3_metas_24_mru <= 1'b0;
        end
        if(_zz_1446) begin
          ways_3_metas_25_mru <= 1'b0;
        end
        if(_zz_1447) begin
          ways_3_metas_26_mru <= 1'b0;
        end
        if(_zz_1448) begin
          ways_3_metas_27_mru <= 1'b0;
        end
        if(_zz_1449) begin
          ways_3_metas_28_mru <= 1'b0;
        end
        if(_zz_1450) begin
          ways_3_metas_29_mru <= 1'b0;
        end
        if(_zz_1451) begin
          ways_3_metas_30_mru <= 1'b0;
        end
        if(_zz_1452) begin
          ways_3_metas_31_mru <= 1'b0;
        end
        if(_zz_1453) begin
          ways_3_metas_32_mru <= 1'b0;
        end
        if(_zz_1454) begin
          ways_3_metas_33_mru <= 1'b0;
        end
        if(_zz_1455) begin
          ways_3_metas_34_mru <= 1'b0;
        end
        if(_zz_1456) begin
          ways_3_metas_35_mru <= 1'b0;
        end
        if(_zz_1457) begin
          ways_3_metas_36_mru <= 1'b0;
        end
        if(_zz_1458) begin
          ways_3_metas_37_mru <= 1'b0;
        end
        if(_zz_1459) begin
          ways_3_metas_38_mru <= 1'b0;
        end
        if(_zz_1460) begin
          ways_3_metas_39_mru <= 1'b0;
        end
        if(_zz_1461) begin
          ways_3_metas_40_mru <= 1'b0;
        end
        if(_zz_1462) begin
          ways_3_metas_41_mru <= 1'b0;
        end
        if(_zz_1463) begin
          ways_3_metas_42_mru <= 1'b0;
        end
        if(_zz_1464) begin
          ways_3_metas_43_mru <= 1'b0;
        end
        if(_zz_1465) begin
          ways_3_metas_44_mru <= 1'b0;
        end
        if(_zz_1466) begin
          ways_3_metas_45_mru <= 1'b0;
        end
        if(_zz_1467) begin
          ways_3_metas_46_mru <= 1'b0;
        end
        if(_zz_1468) begin
          ways_3_metas_47_mru <= 1'b0;
        end
        if(_zz_1469) begin
          ways_3_metas_48_mru <= 1'b0;
        end
        if(_zz_1470) begin
          ways_3_metas_49_mru <= 1'b0;
        end
        if(_zz_1471) begin
          ways_3_metas_50_mru <= 1'b0;
        end
        if(_zz_1472) begin
          ways_3_metas_51_mru <= 1'b0;
        end
        if(_zz_1473) begin
          ways_3_metas_52_mru <= 1'b0;
        end
        if(_zz_1474) begin
          ways_3_metas_53_mru <= 1'b0;
        end
        if(_zz_1475) begin
          ways_3_metas_54_mru <= 1'b0;
        end
        if(_zz_1476) begin
          ways_3_metas_55_mru <= 1'b0;
        end
        if(_zz_1477) begin
          ways_3_metas_56_mru <= 1'b0;
        end
        if(_zz_1478) begin
          ways_3_metas_57_mru <= 1'b0;
        end
        if(_zz_1479) begin
          ways_3_metas_58_mru <= 1'b0;
        end
        if(_zz_1480) begin
          ways_3_metas_59_mru <= 1'b0;
        end
        if(_zz_1481) begin
          ways_3_metas_60_mru <= 1'b0;
        end
        if(_zz_1482) begin
          ways_3_metas_61_mru <= 1'b0;
        end
        if(_zz_1483) begin
          ways_3_metas_62_mru <= 1'b0;
        end
        if(_zz_1484) begin
          ways_3_metas_63_mru <= 1'b0;
        end
        if(_zz_1485) begin
          ways_3_metas_64_mru <= 1'b0;
        end
        if(_zz_1486) begin
          ways_3_metas_65_mru <= 1'b0;
        end
        if(_zz_1487) begin
          ways_3_metas_66_mru <= 1'b0;
        end
        if(_zz_1488) begin
          ways_3_metas_67_mru <= 1'b0;
        end
        if(_zz_1489) begin
          ways_3_metas_68_mru <= 1'b0;
        end
        if(_zz_1490) begin
          ways_3_metas_69_mru <= 1'b0;
        end
        if(_zz_1491) begin
          ways_3_metas_70_mru <= 1'b0;
        end
        if(_zz_1492) begin
          ways_3_metas_71_mru <= 1'b0;
        end
        if(_zz_1493) begin
          ways_3_metas_72_mru <= 1'b0;
        end
        if(_zz_1494) begin
          ways_3_metas_73_mru <= 1'b0;
        end
        if(_zz_1495) begin
          ways_3_metas_74_mru <= 1'b0;
        end
        if(_zz_1496) begin
          ways_3_metas_75_mru <= 1'b0;
        end
        if(_zz_1497) begin
          ways_3_metas_76_mru <= 1'b0;
        end
        if(_zz_1498) begin
          ways_3_metas_77_mru <= 1'b0;
        end
        if(_zz_1499) begin
          ways_3_metas_78_mru <= 1'b0;
        end
        if(_zz_1500) begin
          ways_3_metas_79_mru <= 1'b0;
        end
        if(_zz_1501) begin
          ways_3_metas_80_mru <= 1'b0;
        end
        if(_zz_1502) begin
          ways_3_metas_81_mru <= 1'b0;
        end
        if(_zz_1503) begin
          ways_3_metas_82_mru <= 1'b0;
        end
        if(_zz_1504) begin
          ways_3_metas_83_mru <= 1'b0;
        end
        if(_zz_1505) begin
          ways_3_metas_84_mru <= 1'b0;
        end
        if(_zz_1506) begin
          ways_3_metas_85_mru <= 1'b0;
        end
        if(_zz_1507) begin
          ways_3_metas_86_mru <= 1'b0;
        end
        if(_zz_1508) begin
          ways_3_metas_87_mru <= 1'b0;
        end
        if(_zz_1509) begin
          ways_3_metas_88_mru <= 1'b0;
        end
        if(_zz_1510) begin
          ways_3_metas_89_mru <= 1'b0;
        end
        if(_zz_1511) begin
          ways_3_metas_90_mru <= 1'b0;
        end
        if(_zz_1512) begin
          ways_3_metas_91_mru <= 1'b0;
        end
        if(_zz_1513) begin
          ways_3_metas_92_mru <= 1'b0;
        end
        if(_zz_1514) begin
          ways_3_metas_93_mru <= 1'b0;
        end
        if(_zz_1515) begin
          ways_3_metas_94_mru <= 1'b0;
        end
        if(_zz_1516) begin
          ways_3_metas_95_mru <= 1'b0;
        end
        if(_zz_1517) begin
          ways_3_metas_96_mru <= 1'b0;
        end
        if(_zz_1518) begin
          ways_3_metas_97_mru <= 1'b0;
        end
        if(_zz_1519) begin
          ways_3_metas_98_mru <= 1'b0;
        end
        if(_zz_1520) begin
          ways_3_metas_99_mru <= 1'b0;
        end
        if(_zz_1521) begin
          ways_3_metas_100_mru <= 1'b0;
        end
        if(_zz_1522) begin
          ways_3_metas_101_mru <= 1'b0;
        end
        if(_zz_1523) begin
          ways_3_metas_102_mru <= 1'b0;
        end
        if(_zz_1524) begin
          ways_3_metas_103_mru <= 1'b0;
        end
        if(_zz_1525) begin
          ways_3_metas_104_mru <= 1'b0;
        end
        if(_zz_1526) begin
          ways_3_metas_105_mru <= 1'b0;
        end
        if(_zz_1527) begin
          ways_3_metas_106_mru <= 1'b0;
        end
        if(_zz_1528) begin
          ways_3_metas_107_mru <= 1'b0;
        end
        if(_zz_1529) begin
          ways_3_metas_108_mru <= 1'b0;
        end
        if(_zz_1530) begin
          ways_3_metas_109_mru <= 1'b0;
        end
        if(_zz_1531) begin
          ways_3_metas_110_mru <= 1'b0;
        end
        if(_zz_1532) begin
          ways_3_metas_111_mru <= 1'b0;
        end
        if(_zz_1533) begin
          ways_3_metas_112_mru <= 1'b0;
        end
        if(_zz_1534) begin
          ways_3_metas_113_mru <= 1'b0;
        end
        if(_zz_1535) begin
          ways_3_metas_114_mru <= 1'b0;
        end
        if(_zz_1536) begin
          ways_3_metas_115_mru <= 1'b0;
        end
        if(_zz_1537) begin
          ways_3_metas_116_mru <= 1'b0;
        end
        if(_zz_1538) begin
          ways_3_metas_117_mru <= 1'b0;
        end
        if(_zz_1539) begin
          ways_3_metas_118_mru <= 1'b0;
        end
        if(_zz_1540) begin
          ways_3_metas_119_mru <= 1'b0;
        end
        if(_zz_1541) begin
          ways_3_metas_120_mru <= 1'b0;
        end
        if(_zz_1542) begin
          ways_3_metas_121_mru <= 1'b0;
        end
        if(_zz_1543) begin
          ways_3_metas_122_mru <= 1'b0;
        end
        if(_zz_1544) begin
          ways_3_metas_123_mru <= 1'b0;
        end
        if(_zz_1545) begin
          ways_3_metas_124_mru <= 1'b0;
        end
        if(_zz_1546) begin
          ways_3_metas_125_mru <= 1'b0;
        end
        if(_zz_1547) begin
          ways_3_metas_126_mru <= 1'b0;
        end
        if(_zz_1548) begin
          ways_3_metas_127_mru <= 1'b0;
        end
        if(_zz_1421) begin
          ways_3_metas_0_vld <= 1'b0;
        end
        if(_zz_1422) begin
          ways_3_metas_1_vld <= 1'b0;
        end
        if(_zz_1423) begin
          ways_3_metas_2_vld <= 1'b0;
        end
        if(_zz_1424) begin
          ways_3_metas_3_vld <= 1'b0;
        end
        if(_zz_1425) begin
          ways_3_metas_4_vld <= 1'b0;
        end
        if(_zz_1426) begin
          ways_3_metas_5_vld <= 1'b0;
        end
        if(_zz_1427) begin
          ways_3_metas_6_vld <= 1'b0;
        end
        if(_zz_1428) begin
          ways_3_metas_7_vld <= 1'b0;
        end
        if(_zz_1429) begin
          ways_3_metas_8_vld <= 1'b0;
        end
        if(_zz_1430) begin
          ways_3_metas_9_vld <= 1'b0;
        end
        if(_zz_1431) begin
          ways_3_metas_10_vld <= 1'b0;
        end
        if(_zz_1432) begin
          ways_3_metas_11_vld <= 1'b0;
        end
        if(_zz_1433) begin
          ways_3_metas_12_vld <= 1'b0;
        end
        if(_zz_1434) begin
          ways_3_metas_13_vld <= 1'b0;
        end
        if(_zz_1435) begin
          ways_3_metas_14_vld <= 1'b0;
        end
        if(_zz_1436) begin
          ways_3_metas_15_vld <= 1'b0;
        end
        if(_zz_1437) begin
          ways_3_metas_16_vld <= 1'b0;
        end
        if(_zz_1438) begin
          ways_3_metas_17_vld <= 1'b0;
        end
        if(_zz_1439) begin
          ways_3_metas_18_vld <= 1'b0;
        end
        if(_zz_1440) begin
          ways_3_metas_19_vld <= 1'b0;
        end
        if(_zz_1441) begin
          ways_3_metas_20_vld <= 1'b0;
        end
        if(_zz_1442) begin
          ways_3_metas_21_vld <= 1'b0;
        end
        if(_zz_1443) begin
          ways_3_metas_22_vld <= 1'b0;
        end
        if(_zz_1444) begin
          ways_3_metas_23_vld <= 1'b0;
        end
        if(_zz_1445) begin
          ways_3_metas_24_vld <= 1'b0;
        end
        if(_zz_1446) begin
          ways_3_metas_25_vld <= 1'b0;
        end
        if(_zz_1447) begin
          ways_3_metas_26_vld <= 1'b0;
        end
        if(_zz_1448) begin
          ways_3_metas_27_vld <= 1'b0;
        end
        if(_zz_1449) begin
          ways_3_metas_28_vld <= 1'b0;
        end
        if(_zz_1450) begin
          ways_3_metas_29_vld <= 1'b0;
        end
        if(_zz_1451) begin
          ways_3_metas_30_vld <= 1'b0;
        end
        if(_zz_1452) begin
          ways_3_metas_31_vld <= 1'b0;
        end
        if(_zz_1453) begin
          ways_3_metas_32_vld <= 1'b0;
        end
        if(_zz_1454) begin
          ways_3_metas_33_vld <= 1'b0;
        end
        if(_zz_1455) begin
          ways_3_metas_34_vld <= 1'b0;
        end
        if(_zz_1456) begin
          ways_3_metas_35_vld <= 1'b0;
        end
        if(_zz_1457) begin
          ways_3_metas_36_vld <= 1'b0;
        end
        if(_zz_1458) begin
          ways_3_metas_37_vld <= 1'b0;
        end
        if(_zz_1459) begin
          ways_3_metas_38_vld <= 1'b0;
        end
        if(_zz_1460) begin
          ways_3_metas_39_vld <= 1'b0;
        end
        if(_zz_1461) begin
          ways_3_metas_40_vld <= 1'b0;
        end
        if(_zz_1462) begin
          ways_3_metas_41_vld <= 1'b0;
        end
        if(_zz_1463) begin
          ways_3_metas_42_vld <= 1'b0;
        end
        if(_zz_1464) begin
          ways_3_metas_43_vld <= 1'b0;
        end
        if(_zz_1465) begin
          ways_3_metas_44_vld <= 1'b0;
        end
        if(_zz_1466) begin
          ways_3_metas_45_vld <= 1'b0;
        end
        if(_zz_1467) begin
          ways_3_metas_46_vld <= 1'b0;
        end
        if(_zz_1468) begin
          ways_3_metas_47_vld <= 1'b0;
        end
        if(_zz_1469) begin
          ways_3_metas_48_vld <= 1'b0;
        end
        if(_zz_1470) begin
          ways_3_metas_49_vld <= 1'b0;
        end
        if(_zz_1471) begin
          ways_3_metas_50_vld <= 1'b0;
        end
        if(_zz_1472) begin
          ways_3_metas_51_vld <= 1'b0;
        end
        if(_zz_1473) begin
          ways_3_metas_52_vld <= 1'b0;
        end
        if(_zz_1474) begin
          ways_3_metas_53_vld <= 1'b0;
        end
        if(_zz_1475) begin
          ways_3_metas_54_vld <= 1'b0;
        end
        if(_zz_1476) begin
          ways_3_metas_55_vld <= 1'b0;
        end
        if(_zz_1477) begin
          ways_3_metas_56_vld <= 1'b0;
        end
        if(_zz_1478) begin
          ways_3_metas_57_vld <= 1'b0;
        end
        if(_zz_1479) begin
          ways_3_metas_58_vld <= 1'b0;
        end
        if(_zz_1480) begin
          ways_3_metas_59_vld <= 1'b0;
        end
        if(_zz_1481) begin
          ways_3_metas_60_vld <= 1'b0;
        end
        if(_zz_1482) begin
          ways_3_metas_61_vld <= 1'b0;
        end
        if(_zz_1483) begin
          ways_3_metas_62_vld <= 1'b0;
        end
        if(_zz_1484) begin
          ways_3_metas_63_vld <= 1'b0;
        end
        if(_zz_1485) begin
          ways_3_metas_64_vld <= 1'b0;
        end
        if(_zz_1486) begin
          ways_3_metas_65_vld <= 1'b0;
        end
        if(_zz_1487) begin
          ways_3_metas_66_vld <= 1'b0;
        end
        if(_zz_1488) begin
          ways_3_metas_67_vld <= 1'b0;
        end
        if(_zz_1489) begin
          ways_3_metas_68_vld <= 1'b0;
        end
        if(_zz_1490) begin
          ways_3_metas_69_vld <= 1'b0;
        end
        if(_zz_1491) begin
          ways_3_metas_70_vld <= 1'b0;
        end
        if(_zz_1492) begin
          ways_3_metas_71_vld <= 1'b0;
        end
        if(_zz_1493) begin
          ways_3_metas_72_vld <= 1'b0;
        end
        if(_zz_1494) begin
          ways_3_metas_73_vld <= 1'b0;
        end
        if(_zz_1495) begin
          ways_3_metas_74_vld <= 1'b0;
        end
        if(_zz_1496) begin
          ways_3_metas_75_vld <= 1'b0;
        end
        if(_zz_1497) begin
          ways_3_metas_76_vld <= 1'b0;
        end
        if(_zz_1498) begin
          ways_3_metas_77_vld <= 1'b0;
        end
        if(_zz_1499) begin
          ways_3_metas_78_vld <= 1'b0;
        end
        if(_zz_1500) begin
          ways_3_metas_79_vld <= 1'b0;
        end
        if(_zz_1501) begin
          ways_3_metas_80_vld <= 1'b0;
        end
        if(_zz_1502) begin
          ways_3_metas_81_vld <= 1'b0;
        end
        if(_zz_1503) begin
          ways_3_metas_82_vld <= 1'b0;
        end
        if(_zz_1504) begin
          ways_3_metas_83_vld <= 1'b0;
        end
        if(_zz_1505) begin
          ways_3_metas_84_vld <= 1'b0;
        end
        if(_zz_1506) begin
          ways_3_metas_85_vld <= 1'b0;
        end
        if(_zz_1507) begin
          ways_3_metas_86_vld <= 1'b0;
        end
        if(_zz_1508) begin
          ways_3_metas_87_vld <= 1'b0;
        end
        if(_zz_1509) begin
          ways_3_metas_88_vld <= 1'b0;
        end
        if(_zz_1510) begin
          ways_3_metas_89_vld <= 1'b0;
        end
        if(_zz_1511) begin
          ways_3_metas_90_vld <= 1'b0;
        end
        if(_zz_1512) begin
          ways_3_metas_91_vld <= 1'b0;
        end
        if(_zz_1513) begin
          ways_3_metas_92_vld <= 1'b0;
        end
        if(_zz_1514) begin
          ways_3_metas_93_vld <= 1'b0;
        end
        if(_zz_1515) begin
          ways_3_metas_94_vld <= 1'b0;
        end
        if(_zz_1516) begin
          ways_3_metas_95_vld <= 1'b0;
        end
        if(_zz_1517) begin
          ways_3_metas_96_vld <= 1'b0;
        end
        if(_zz_1518) begin
          ways_3_metas_97_vld <= 1'b0;
        end
        if(_zz_1519) begin
          ways_3_metas_98_vld <= 1'b0;
        end
        if(_zz_1520) begin
          ways_3_metas_99_vld <= 1'b0;
        end
        if(_zz_1521) begin
          ways_3_metas_100_vld <= 1'b0;
        end
        if(_zz_1522) begin
          ways_3_metas_101_vld <= 1'b0;
        end
        if(_zz_1523) begin
          ways_3_metas_102_vld <= 1'b0;
        end
        if(_zz_1524) begin
          ways_3_metas_103_vld <= 1'b0;
        end
        if(_zz_1525) begin
          ways_3_metas_104_vld <= 1'b0;
        end
        if(_zz_1526) begin
          ways_3_metas_105_vld <= 1'b0;
        end
        if(_zz_1527) begin
          ways_3_metas_106_vld <= 1'b0;
        end
        if(_zz_1528) begin
          ways_3_metas_107_vld <= 1'b0;
        end
        if(_zz_1529) begin
          ways_3_metas_108_vld <= 1'b0;
        end
        if(_zz_1530) begin
          ways_3_metas_109_vld <= 1'b0;
        end
        if(_zz_1531) begin
          ways_3_metas_110_vld <= 1'b0;
        end
        if(_zz_1532) begin
          ways_3_metas_111_vld <= 1'b0;
        end
        if(_zz_1533) begin
          ways_3_metas_112_vld <= 1'b0;
        end
        if(_zz_1534) begin
          ways_3_metas_113_vld <= 1'b0;
        end
        if(_zz_1535) begin
          ways_3_metas_114_vld <= 1'b0;
        end
        if(_zz_1536) begin
          ways_3_metas_115_vld <= 1'b0;
        end
        if(_zz_1537) begin
          ways_3_metas_116_vld <= 1'b0;
        end
        if(_zz_1538) begin
          ways_3_metas_117_vld <= 1'b0;
        end
        if(_zz_1539) begin
          ways_3_metas_118_vld <= 1'b0;
        end
        if(_zz_1540) begin
          ways_3_metas_119_vld <= 1'b0;
        end
        if(_zz_1541) begin
          ways_3_metas_120_vld <= 1'b0;
        end
        if(_zz_1542) begin
          ways_3_metas_121_vld <= 1'b0;
        end
        if(_zz_1543) begin
          ways_3_metas_122_vld <= 1'b0;
        end
        if(_zz_1544) begin
          ways_3_metas_123_vld <= 1'b0;
        end
        if(_zz_1545) begin
          ways_3_metas_124_vld <= 1'b0;
        end
        if(_zz_1546) begin
          ways_3_metas_125_vld <= 1'b0;
        end
        if(_zz_1547) begin
          ways_3_metas_126_vld <= 1'b0;
        end
        if(_zz_1548) begin
          ways_3_metas_127_vld <= 1'b0;
        end
      end else begin
        if(when_ICache_l210_3) begin
          if(cache_hit_3) begin
            if(_zz_1163) begin
              ways_3_metas_0_mru <= 1'b1;
            end
            if(_zz_1164) begin
              ways_3_metas_1_mru <= 1'b1;
            end
            if(_zz_1165) begin
              ways_3_metas_2_mru <= 1'b1;
            end
            if(_zz_1166) begin
              ways_3_metas_3_mru <= 1'b1;
            end
            if(_zz_1167) begin
              ways_3_metas_4_mru <= 1'b1;
            end
            if(_zz_1168) begin
              ways_3_metas_5_mru <= 1'b1;
            end
            if(_zz_1169) begin
              ways_3_metas_6_mru <= 1'b1;
            end
            if(_zz_1170) begin
              ways_3_metas_7_mru <= 1'b1;
            end
            if(_zz_1171) begin
              ways_3_metas_8_mru <= 1'b1;
            end
            if(_zz_1172) begin
              ways_3_metas_9_mru <= 1'b1;
            end
            if(_zz_1173) begin
              ways_3_metas_10_mru <= 1'b1;
            end
            if(_zz_1174) begin
              ways_3_metas_11_mru <= 1'b1;
            end
            if(_zz_1175) begin
              ways_3_metas_12_mru <= 1'b1;
            end
            if(_zz_1176) begin
              ways_3_metas_13_mru <= 1'b1;
            end
            if(_zz_1177) begin
              ways_3_metas_14_mru <= 1'b1;
            end
            if(_zz_1178) begin
              ways_3_metas_15_mru <= 1'b1;
            end
            if(_zz_1179) begin
              ways_3_metas_16_mru <= 1'b1;
            end
            if(_zz_1180) begin
              ways_3_metas_17_mru <= 1'b1;
            end
            if(_zz_1181) begin
              ways_3_metas_18_mru <= 1'b1;
            end
            if(_zz_1182) begin
              ways_3_metas_19_mru <= 1'b1;
            end
            if(_zz_1183) begin
              ways_3_metas_20_mru <= 1'b1;
            end
            if(_zz_1184) begin
              ways_3_metas_21_mru <= 1'b1;
            end
            if(_zz_1185) begin
              ways_3_metas_22_mru <= 1'b1;
            end
            if(_zz_1186) begin
              ways_3_metas_23_mru <= 1'b1;
            end
            if(_zz_1187) begin
              ways_3_metas_24_mru <= 1'b1;
            end
            if(_zz_1188) begin
              ways_3_metas_25_mru <= 1'b1;
            end
            if(_zz_1189) begin
              ways_3_metas_26_mru <= 1'b1;
            end
            if(_zz_1190) begin
              ways_3_metas_27_mru <= 1'b1;
            end
            if(_zz_1191) begin
              ways_3_metas_28_mru <= 1'b1;
            end
            if(_zz_1192) begin
              ways_3_metas_29_mru <= 1'b1;
            end
            if(_zz_1193) begin
              ways_3_metas_30_mru <= 1'b1;
            end
            if(_zz_1194) begin
              ways_3_metas_31_mru <= 1'b1;
            end
            if(_zz_1195) begin
              ways_3_metas_32_mru <= 1'b1;
            end
            if(_zz_1196) begin
              ways_3_metas_33_mru <= 1'b1;
            end
            if(_zz_1197) begin
              ways_3_metas_34_mru <= 1'b1;
            end
            if(_zz_1198) begin
              ways_3_metas_35_mru <= 1'b1;
            end
            if(_zz_1199) begin
              ways_3_metas_36_mru <= 1'b1;
            end
            if(_zz_1200) begin
              ways_3_metas_37_mru <= 1'b1;
            end
            if(_zz_1201) begin
              ways_3_metas_38_mru <= 1'b1;
            end
            if(_zz_1202) begin
              ways_3_metas_39_mru <= 1'b1;
            end
            if(_zz_1203) begin
              ways_3_metas_40_mru <= 1'b1;
            end
            if(_zz_1204) begin
              ways_3_metas_41_mru <= 1'b1;
            end
            if(_zz_1205) begin
              ways_3_metas_42_mru <= 1'b1;
            end
            if(_zz_1206) begin
              ways_3_metas_43_mru <= 1'b1;
            end
            if(_zz_1207) begin
              ways_3_metas_44_mru <= 1'b1;
            end
            if(_zz_1208) begin
              ways_3_metas_45_mru <= 1'b1;
            end
            if(_zz_1209) begin
              ways_3_metas_46_mru <= 1'b1;
            end
            if(_zz_1210) begin
              ways_3_metas_47_mru <= 1'b1;
            end
            if(_zz_1211) begin
              ways_3_metas_48_mru <= 1'b1;
            end
            if(_zz_1212) begin
              ways_3_metas_49_mru <= 1'b1;
            end
            if(_zz_1213) begin
              ways_3_metas_50_mru <= 1'b1;
            end
            if(_zz_1214) begin
              ways_3_metas_51_mru <= 1'b1;
            end
            if(_zz_1215) begin
              ways_3_metas_52_mru <= 1'b1;
            end
            if(_zz_1216) begin
              ways_3_metas_53_mru <= 1'b1;
            end
            if(_zz_1217) begin
              ways_3_metas_54_mru <= 1'b1;
            end
            if(_zz_1218) begin
              ways_3_metas_55_mru <= 1'b1;
            end
            if(_zz_1219) begin
              ways_3_metas_56_mru <= 1'b1;
            end
            if(_zz_1220) begin
              ways_3_metas_57_mru <= 1'b1;
            end
            if(_zz_1221) begin
              ways_3_metas_58_mru <= 1'b1;
            end
            if(_zz_1222) begin
              ways_3_metas_59_mru <= 1'b1;
            end
            if(_zz_1223) begin
              ways_3_metas_60_mru <= 1'b1;
            end
            if(_zz_1224) begin
              ways_3_metas_61_mru <= 1'b1;
            end
            if(_zz_1225) begin
              ways_3_metas_62_mru <= 1'b1;
            end
            if(_zz_1226) begin
              ways_3_metas_63_mru <= 1'b1;
            end
            if(_zz_1227) begin
              ways_3_metas_64_mru <= 1'b1;
            end
            if(_zz_1228) begin
              ways_3_metas_65_mru <= 1'b1;
            end
            if(_zz_1229) begin
              ways_3_metas_66_mru <= 1'b1;
            end
            if(_zz_1230) begin
              ways_3_metas_67_mru <= 1'b1;
            end
            if(_zz_1231) begin
              ways_3_metas_68_mru <= 1'b1;
            end
            if(_zz_1232) begin
              ways_3_metas_69_mru <= 1'b1;
            end
            if(_zz_1233) begin
              ways_3_metas_70_mru <= 1'b1;
            end
            if(_zz_1234) begin
              ways_3_metas_71_mru <= 1'b1;
            end
            if(_zz_1235) begin
              ways_3_metas_72_mru <= 1'b1;
            end
            if(_zz_1236) begin
              ways_3_metas_73_mru <= 1'b1;
            end
            if(_zz_1237) begin
              ways_3_metas_74_mru <= 1'b1;
            end
            if(_zz_1238) begin
              ways_3_metas_75_mru <= 1'b1;
            end
            if(_zz_1239) begin
              ways_3_metas_76_mru <= 1'b1;
            end
            if(_zz_1240) begin
              ways_3_metas_77_mru <= 1'b1;
            end
            if(_zz_1241) begin
              ways_3_metas_78_mru <= 1'b1;
            end
            if(_zz_1242) begin
              ways_3_metas_79_mru <= 1'b1;
            end
            if(_zz_1243) begin
              ways_3_metas_80_mru <= 1'b1;
            end
            if(_zz_1244) begin
              ways_3_metas_81_mru <= 1'b1;
            end
            if(_zz_1245) begin
              ways_3_metas_82_mru <= 1'b1;
            end
            if(_zz_1246) begin
              ways_3_metas_83_mru <= 1'b1;
            end
            if(_zz_1247) begin
              ways_3_metas_84_mru <= 1'b1;
            end
            if(_zz_1248) begin
              ways_3_metas_85_mru <= 1'b1;
            end
            if(_zz_1249) begin
              ways_3_metas_86_mru <= 1'b1;
            end
            if(_zz_1250) begin
              ways_3_metas_87_mru <= 1'b1;
            end
            if(_zz_1251) begin
              ways_3_metas_88_mru <= 1'b1;
            end
            if(_zz_1252) begin
              ways_3_metas_89_mru <= 1'b1;
            end
            if(_zz_1253) begin
              ways_3_metas_90_mru <= 1'b1;
            end
            if(_zz_1254) begin
              ways_3_metas_91_mru <= 1'b1;
            end
            if(_zz_1255) begin
              ways_3_metas_92_mru <= 1'b1;
            end
            if(_zz_1256) begin
              ways_3_metas_93_mru <= 1'b1;
            end
            if(_zz_1257) begin
              ways_3_metas_94_mru <= 1'b1;
            end
            if(_zz_1258) begin
              ways_3_metas_95_mru <= 1'b1;
            end
            if(_zz_1259) begin
              ways_3_metas_96_mru <= 1'b1;
            end
            if(_zz_1260) begin
              ways_3_metas_97_mru <= 1'b1;
            end
            if(_zz_1261) begin
              ways_3_metas_98_mru <= 1'b1;
            end
            if(_zz_1262) begin
              ways_3_metas_99_mru <= 1'b1;
            end
            if(_zz_1263) begin
              ways_3_metas_100_mru <= 1'b1;
            end
            if(_zz_1264) begin
              ways_3_metas_101_mru <= 1'b1;
            end
            if(_zz_1265) begin
              ways_3_metas_102_mru <= 1'b1;
            end
            if(_zz_1266) begin
              ways_3_metas_103_mru <= 1'b1;
            end
            if(_zz_1267) begin
              ways_3_metas_104_mru <= 1'b1;
            end
            if(_zz_1268) begin
              ways_3_metas_105_mru <= 1'b1;
            end
            if(_zz_1269) begin
              ways_3_metas_106_mru <= 1'b1;
            end
            if(_zz_1270) begin
              ways_3_metas_107_mru <= 1'b1;
            end
            if(_zz_1271) begin
              ways_3_metas_108_mru <= 1'b1;
            end
            if(_zz_1272) begin
              ways_3_metas_109_mru <= 1'b1;
            end
            if(_zz_1273) begin
              ways_3_metas_110_mru <= 1'b1;
            end
            if(_zz_1274) begin
              ways_3_metas_111_mru <= 1'b1;
            end
            if(_zz_1275) begin
              ways_3_metas_112_mru <= 1'b1;
            end
            if(_zz_1276) begin
              ways_3_metas_113_mru <= 1'b1;
            end
            if(_zz_1277) begin
              ways_3_metas_114_mru <= 1'b1;
            end
            if(_zz_1278) begin
              ways_3_metas_115_mru <= 1'b1;
            end
            if(_zz_1279) begin
              ways_3_metas_116_mru <= 1'b1;
            end
            if(_zz_1280) begin
              ways_3_metas_117_mru <= 1'b1;
            end
            if(_zz_1281) begin
              ways_3_metas_118_mru <= 1'b1;
            end
            if(_zz_1282) begin
              ways_3_metas_119_mru <= 1'b1;
            end
            if(_zz_1283) begin
              ways_3_metas_120_mru <= 1'b1;
            end
            if(_zz_1284) begin
              ways_3_metas_121_mru <= 1'b1;
            end
            if(_zz_1285) begin
              ways_3_metas_122_mru <= 1'b1;
            end
            if(_zz_1286) begin
              ways_3_metas_123_mru <= 1'b1;
            end
            if(_zz_1287) begin
              ways_3_metas_124_mru <= 1'b1;
            end
            if(_zz_1288) begin
              ways_3_metas_125_mru <= 1'b1;
            end
            if(_zz_1289) begin
              ways_3_metas_126_mru <= 1'b1;
            end
            if(_zz_1290) begin
              ways_3_metas_127_mru <= 1'b1;
            end
          end else begin
            if(_zz_1163) begin
              ways_3_metas_0_mru <= 1'b0;
            end
            if(_zz_1164) begin
              ways_3_metas_1_mru <= 1'b0;
            end
            if(_zz_1165) begin
              ways_3_metas_2_mru <= 1'b0;
            end
            if(_zz_1166) begin
              ways_3_metas_3_mru <= 1'b0;
            end
            if(_zz_1167) begin
              ways_3_metas_4_mru <= 1'b0;
            end
            if(_zz_1168) begin
              ways_3_metas_5_mru <= 1'b0;
            end
            if(_zz_1169) begin
              ways_3_metas_6_mru <= 1'b0;
            end
            if(_zz_1170) begin
              ways_3_metas_7_mru <= 1'b0;
            end
            if(_zz_1171) begin
              ways_3_metas_8_mru <= 1'b0;
            end
            if(_zz_1172) begin
              ways_3_metas_9_mru <= 1'b0;
            end
            if(_zz_1173) begin
              ways_3_metas_10_mru <= 1'b0;
            end
            if(_zz_1174) begin
              ways_3_metas_11_mru <= 1'b0;
            end
            if(_zz_1175) begin
              ways_3_metas_12_mru <= 1'b0;
            end
            if(_zz_1176) begin
              ways_3_metas_13_mru <= 1'b0;
            end
            if(_zz_1177) begin
              ways_3_metas_14_mru <= 1'b0;
            end
            if(_zz_1178) begin
              ways_3_metas_15_mru <= 1'b0;
            end
            if(_zz_1179) begin
              ways_3_metas_16_mru <= 1'b0;
            end
            if(_zz_1180) begin
              ways_3_metas_17_mru <= 1'b0;
            end
            if(_zz_1181) begin
              ways_3_metas_18_mru <= 1'b0;
            end
            if(_zz_1182) begin
              ways_3_metas_19_mru <= 1'b0;
            end
            if(_zz_1183) begin
              ways_3_metas_20_mru <= 1'b0;
            end
            if(_zz_1184) begin
              ways_3_metas_21_mru <= 1'b0;
            end
            if(_zz_1185) begin
              ways_3_metas_22_mru <= 1'b0;
            end
            if(_zz_1186) begin
              ways_3_metas_23_mru <= 1'b0;
            end
            if(_zz_1187) begin
              ways_3_metas_24_mru <= 1'b0;
            end
            if(_zz_1188) begin
              ways_3_metas_25_mru <= 1'b0;
            end
            if(_zz_1189) begin
              ways_3_metas_26_mru <= 1'b0;
            end
            if(_zz_1190) begin
              ways_3_metas_27_mru <= 1'b0;
            end
            if(_zz_1191) begin
              ways_3_metas_28_mru <= 1'b0;
            end
            if(_zz_1192) begin
              ways_3_metas_29_mru <= 1'b0;
            end
            if(_zz_1193) begin
              ways_3_metas_30_mru <= 1'b0;
            end
            if(_zz_1194) begin
              ways_3_metas_31_mru <= 1'b0;
            end
            if(_zz_1195) begin
              ways_3_metas_32_mru <= 1'b0;
            end
            if(_zz_1196) begin
              ways_3_metas_33_mru <= 1'b0;
            end
            if(_zz_1197) begin
              ways_3_metas_34_mru <= 1'b0;
            end
            if(_zz_1198) begin
              ways_3_metas_35_mru <= 1'b0;
            end
            if(_zz_1199) begin
              ways_3_metas_36_mru <= 1'b0;
            end
            if(_zz_1200) begin
              ways_3_metas_37_mru <= 1'b0;
            end
            if(_zz_1201) begin
              ways_3_metas_38_mru <= 1'b0;
            end
            if(_zz_1202) begin
              ways_3_metas_39_mru <= 1'b0;
            end
            if(_zz_1203) begin
              ways_3_metas_40_mru <= 1'b0;
            end
            if(_zz_1204) begin
              ways_3_metas_41_mru <= 1'b0;
            end
            if(_zz_1205) begin
              ways_3_metas_42_mru <= 1'b0;
            end
            if(_zz_1206) begin
              ways_3_metas_43_mru <= 1'b0;
            end
            if(_zz_1207) begin
              ways_3_metas_44_mru <= 1'b0;
            end
            if(_zz_1208) begin
              ways_3_metas_45_mru <= 1'b0;
            end
            if(_zz_1209) begin
              ways_3_metas_46_mru <= 1'b0;
            end
            if(_zz_1210) begin
              ways_3_metas_47_mru <= 1'b0;
            end
            if(_zz_1211) begin
              ways_3_metas_48_mru <= 1'b0;
            end
            if(_zz_1212) begin
              ways_3_metas_49_mru <= 1'b0;
            end
            if(_zz_1213) begin
              ways_3_metas_50_mru <= 1'b0;
            end
            if(_zz_1214) begin
              ways_3_metas_51_mru <= 1'b0;
            end
            if(_zz_1215) begin
              ways_3_metas_52_mru <= 1'b0;
            end
            if(_zz_1216) begin
              ways_3_metas_53_mru <= 1'b0;
            end
            if(_zz_1217) begin
              ways_3_metas_54_mru <= 1'b0;
            end
            if(_zz_1218) begin
              ways_3_metas_55_mru <= 1'b0;
            end
            if(_zz_1219) begin
              ways_3_metas_56_mru <= 1'b0;
            end
            if(_zz_1220) begin
              ways_3_metas_57_mru <= 1'b0;
            end
            if(_zz_1221) begin
              ways_3_metas_58_mru <= 1'b0;
            end
            if(_zz_1222) begin
              ways_3_metas_59_mru <= 1'b0;
            end
            if(_zz_1223) begin
              ways_3_metas_60_mru <= 1'b0;
            end
            if(_zz_1224) begin
              ways_3_metas_61_mru <= 1'b0;
            end
            if(_zz_1225) begin
              ways_3_metas_62_mru <= 1'b0;
            end
            if(_zz_1226) begin
              ways_3_metas_63_mru <= 1'b0;
            end
            if(_zz_1227) begin
              ways_3_metas_64_mru <= 1'b0;
            end
            if(_zz_1228) begin
              ways_3_metas_65_mru <= 1'b0;
            end
            if(_zz_1229) begin
              ways_3_metas_66_mru <= 1'b0;
            end
            if(_zz_1230) begin
              ways_3_metas_67_mru <= 1'b0;
            end
            if(_zz_1231) begin
              ways_3_metas_68_mru <= 1'b0;
            end
            if(_zz_1232) begin
              ways_3_metas_69_mru <= 1'b0;
            end
            if(_zz_1233) begin
              ways_3_metas_70_mru <= 1'b0;
            end
            if(_zz_1234) begin
              ways_3_metas_71_mru <= 1'b0;
            end
            if(_zz_1235) begin
              ways_3_metas_72_mru <= 1'b0;
            end
            if(_zz_1236) begin
              ways_3_metas_73_mru <= 1'b0;
            end
            if(_zz_1237) begin
              ways_3_metas_74_mru <= 1'b0;
            end
            if(_zz_1238) begin
              ways_3_metas_75_mru <= 1'b0;
            end
            if(_zz_1239) begin
              ways_3_metas_76_mru <= 1'b0;
            end
            if(_zz_1240) begin
              ways_3_metas_77_mru <= 1'b0;
            end
            if(_zz_1241) begin
              ways_3_metas_78_mru <= 1'b0;
            end
            if(_zz_1242) begin
              ways_3_metas_79_mru <= 1'b0;
            end
            if(_zz_1243) begin
              ways_3_metas_80_mru <= 1'b0;
            end
            if(_zz_1244) begin
              ways_3_metas_81_mru <= 1'b0;
            end
            if(_zz_1245) begin
              ways_3_metas_82_mru <= 1'b0;
            end
            if(_zz_1246) begin
              ways_3_metas_83_mru <= 1'b0;
            end
            if(_zz_1247) begin
              ways_3_metas_84_mru <= 1'b0;
            end
            if(_zz_1248) begin
              ways_3_metas_85_mru <= 1'b0;
            end
            if(_zz_1249) begin
              ways_3_metas_86_mru <= 1'b0;
            end
            if(_zz_1250) begin
              ways_3_metas_87_mru <= 1'b0;
            end
            if(_zz_1251) begin
              ways_3_metas_88_mru <= 1'b0;
            end
            if(_zz_1252) begin
              ways_3_metas_89_mru <= 1'b0;
            end
            if(_zz_1253) begin
              ways_3_metas_90_mru <= 1'b0;
            end
            if(_zz_1254) begin
              ways_3_metas_91_mru <= 1'b0;
            end
            if(_zz_1255) begin
              ways_3_metas_92_mru <= 1'b0;
            end
            if(_zz_1256) begin
              ways_3_metas_93_mru <= 1'b0;
            end
            if(_zz_1257) begin
              ways_3_metas_94_mru <= 1'b0;
            end
            if(_zz_1258) begin
              ways_3_metas_95_mru <= 1'b0;
            end
            if(_zz_1259) begin
              ways_3_metas_96_mru <= 1'b0;
            end
            if(_zz_1260) begin
              ways_3_metas_97_mru <= 1'b0;
            end
            if(_zz_1261) begin
              ways_3_metas_98_mru <= 1'b0;
            end
            if(_zz_1262) begin
              ways_3_metas_99_mru <= 1'b0;
            end
            if(_zz_1263) begin
              ways_3_metas_100_mru <= 1'b0;
            end
            if(_zz_1264) begin
              ways_3_metas_101_mru <= 1'b0;
            end
            if(_zz_1265) begin
              ways_3_metas_102_mru <= 1'b0;
            end
            if(_zz_1266) begin
              ways_3_metas_103_mru <= 1'b0;
            end
            if(_zz_1267) begin
              ways_3_metas_104_mru <= 1'b0;
            end
            if(_zz_1268) begin
              ways_3_metas_105_mru <= 1'b0;
            end
            if(_zz_1269) begin
              ways_3_metas_106_mru <= 1'b0;
            end
            if(_zz_1270) begin
              ways_3_metas_107_mru <= 1'b0;
            end
            if(_zz_1271) begin
              ways_3_metas_108_mru <= 1'b0;
            end
            if(_zz_1272) begin
              ways_3_metas_109_mru <= 1'b0;
            end
            if(_zz_1273) begin
              ways_3_metas_110_mru <= 1'b0;
            end
            if(_zz_1274) begin
              ways_3_metas_111_mru <= 1'b0;
            end
            if(_zz_1275) begin
              ways_3_metas_112_mru <= 1'b0;
            end
            if(_zz_1276) begin
              ways_3_metas_113_mru <= 1'b0;
            end
            if(_zz_1277) begin
              ways_3_metas_114_mru <= 1'b0;
            end
            if(_zz_1278) begin
              ways_3_metas_115_mru <= 1'b0;
            end
            if(_zz_1279) begin
              ways_3_metas_116_mru <= 1'b0;
            end
            if(_zz_1280) begin
              ways_3_metas_117_mru <= 1'b0;
            end
            if(_zz_1281) begin
              ways_3_metas_118_mru <= 1'b0;
            end
            if(_zz_1282) begin
              ways_3_metas_119_mru <= 1'b0;
            end
            if(_zz_1283) begin
              ways_3_metas_120_mru <= 1'b0;
            end
            if(_zz_1284) begin
              ways_3_metas_121_mru <= 1'b0;
            end
            if(_zz_1285) begin
              ways_3_metas_122_mru <= 1'b0;
            end
            if(_zz_1286) begin
              ways_3_metas_123_mru <= 1'b0;
            end
            if(_zz_1287) begin
              ways_3_metas_124_mru <= 1'b0;
            end
            if(_zz_1288) begin
              ways_3_metas_125_mru <= 1'b0;
            end
            if(_zz_1289) begin
              ways_3_metas_126_mru <= 1'b0;
            end
            if(_zz_1290) begin
              ways_3_metas_127_mru <= 1'b0;
            end
          end
        end else begin
          if(when_ICache_l217_3) begin
            if(_zz_1163) begin
              ways_3_metas_0_mru <= 1'b1;
            end
            if(_zz_1164) begin
              ways_3_metas_1_mru <= 1'b1;
            end
            if(_zz_1165) begin
              ways_3_metas_2_mru <= 1'b1;
            end
            if(_zz_1166) begin
              ways_3_metas_3_mru <= 1'b1;
            end
            if(_zz_1167) begin
              ways_3_metas_4_mru <= 1'b1;
            end
            if(_zz_1168) begin
              ways_3_metas_5_mru <= 1'b1;
            end
            if(_zz_1169) begin
              ways_3_metas_6_mru <= 1'b1;
            end
            if(_zz_1170) begin
              ways_3_metas_7_mru <= 1'b1;
            end
            if(_zz_1171) begin
              ways_3_metas_8_mru <= 1'b1;
            end
            if(_zz_1172) begin
              ways_3_metas_9_mru <= 1'b1;
            end
            if(_zz_1173) begin
              ways_3_metas_10_mru <= 1'b1;
            end
            if(_zz_1174) begin
              ways_3_metas_11_mru <= 1'b1;
            end
            if(_zz_1175) begin
              ways_3_metas_12_mru <= 1'b1;
            end
            if(_zz_1176) begin
              ways_3_metas_13_mru <= 1'b1;
            end
            if(_zz_1177) begin
              ways_3_metas_14_mru <= 1'b1;
            end
            if(_zz_1178) begin
              ways_3_metas_15_mru <= 1'b1;
            end
            if(_zz_1179) begin
              ways_3_metas_16_mru <= 1'b1;
            end
            if(_zz_1180) begin
              ways_3_metas_17_mru <= 1'b1;
            end
            if(_zz_1181) begin
              ways_3_metas_18_mru <= 1'b1;
            end
            if(_zz_1182) begin
              ways_3_metas_19_mru <= 1'b1;
            end
            if(_zz_1183) begin
              ways_3_metas_20_mru <= 1'b1;
            end
            if(_zz_1184) begin
              ways_3_metas_21_mru <= 1'b1;
            end
            if(_zz_1185) begin
              ways_3_metas_22_mru <= 1'b1;
            end
            if(_zz_1186) begin
              ways_3_metas_23_mru <= 1'b1;
            end
            if(_zz_1187) begin
              ways_3_metas_24_mru <= 1'b1;
            end
            if(_zz_1188) begin
              ways_3_metas_25_mru <= 1'b1;
            end
            if(_zz_1189) begin
              ways_3_metas_26_mru <= 1'b1;
            end
            if(_zz_1190) begin
              ways_3_metas_27_mru <= 1'b1;
            end
            if(_zz_1191) begin
              ways_3_metas_28_mru <= 1'b1;
            end
            if(_zz_1192) begin
              ways_3_metas_29_mru <= 1'b1;
            end
            if(_zz_1193) begin
              ways_3_metas_30_mru <= 1'b1;
            end
            if(_zz_1194) begin
              ways_3_metas_31_mru <= 1'b1;
            end
            if(_zz_1195) begin
              ways_3_metas_32_mru <= 1'b1;
            end
            if(_zz_1196) begin
              ways_3_metas_33_mru <= 1'b1;
            end
            if(_zz_1197) begin
              ways_3_metas_34_mru <= 1'b1;
            end
            if(_zz_1198) begin
              ways_3_metas_35_mru <= 1'b1;
            end
            if(_zz_1199) begin
              ways_3_metas_36_mru <= 1'b1;
            end
            if(_zz_1200) begin
              ways_3_metas_37_mru <= 1'b1;
            end
            if(_zz_1201) begin
              ways_3_metas_38_mru <= 1'b1;
            end
            if(_zz_1202) begin
              ways_3_metas_39_mru <= 1'b1;
            end
            if(_zz_1203) begin
              ways_3_metas_40_mru <= 1'b1;
            end
            if(_zz_1204) begin
              ways_3_metas_41_mru <= 1'b1;
            end
            if(_zz_1205) begin
              ways_3_metas_42_mru <= 1'b1;
            end
            if(_zz_1206) begin
              ways_3_metas_43_mru <= 1'b1;
            end
            if(_zz_1207) begin
              ways_3_metas_44_mru <= 1'b1;
            end
            if(_zz_1208) begin
              ways_3_metas_45_mru <= 1'b1;
            end
            if(_zz_1209) begin
              ways_3_metas_46_mru <= 1'b1;
            end
            if(_zz_1210) begin
              ways_3_metas_47_mru <= 1'b1;
            end
            if(_zz_1211) begin
              ways_3_metas_48_mru <= 1'b1;
            end
            if(_zz_1212) begin
              ways_3_metas_49_mru <= 1'b1;
            end
            if(_zz_1213) begin
              ways_3_metas_50_mru <= 1'b1;
            end
            if(_zz_1214) begin
              ways_3_metas_51_mru <= 1'b1;
            end
            if(_zz_1215) begin
              ways_3_metas_52_mru <= 1'b1;
            end
            if(_zz_1216) begin
              ways_3_metas_53_mru <= 1'b1;
            end
            if(_zz_1217) begin
              ways_3_metas_54_mru <= 1'b1;
            end
            if(_zz_1218) begin
              ways_3_metas_55_mru <= 1'b1;
            end
            if(_zz_1219) begin
              ways_3_metas_56_mru <= 1'b1;
            end
            if(_zz_1220) begin
              ways_3_metas_57_mru <= 1'b1;
            end
            if(_zz_1221) begin
              ways_3_metas_58_mru <= 1'b1;
            end
            if(_zz_1222) begin
              ways_3_metas_59_mru <= 1'b1;
            end
            if(_zz_1223) begin
              ways_3_metas_60_mru <= 1'b1;
            end
            if(_zz_1224) begin
              ways_3_metas_61_mru <= 1'b1;
            end
            if(_zz_1225) begin
              ways_3_metas_62_mru <= 1'b1;
            end
            if(_zz_1226) begin
              ways_3_metas_63_mru <= 1'b1;
            end
            if(_zz_1227) begin
              ways_3_metas_64_mru <= 1'b1;
            end
            if(_zz_1228) begin
              ways_3_metas_65_mru <= 1'b1;
            end
            if(_zz_1229) begin
              ways_3_metas_66_mru <= 1'b1;
            end
            if(_zz_1230) begin
              ways_3_metas_67_mru <= 1'b1;
            end
            if(_zz_1231) begin
              ways_3_metas_68_mru <= 1'b1;
            end
            if(_zz_1232) begin
              ways_3_metas_69_mru <= 1'b1;
            end
            if(_zz_1233) begin
              ways_3_metas_70_mru <= 1'b1;
            end
            if(_zz_1234) begin
              ways_3_metas_71_mru <= 1'b1;
            end
            if(_zz_1235) begin
              ways_3_metas_72_mru <= 1'b1;
            end
            if(_zz_1236) begin
              ways_3_metas_73_mru <= 1'b1;
            end
            if(_zz_1237) begin
              ways_3_metas_74_mru <= 1'b1;
            end
            if(_zz_1238) begin
              ways_3_metas_75_mru <= 1'b1;
            end
            if(_zz_1239) begin
              ways_3_metas_76_mru <= 1'b1;
            end
            if(_zz_1240) begin
              ways_3_metas_77_mru <= 1'b1;
            end
            if(_zz_1241) begin
              ways_3_metas_78_mru <= 1'b1;
            end
            if(_zz_1242) begin
              ways_3_metas_79_mru <= 1'b1;
            end
            if(_zz_1243) begin
              ways_3_metas_80_mru <= 1'b1;
            end
            if(_zz_1244) begin
              ways_3_metas_81_mru <= 1'b1;
            end
            if(_zz_1245) begin
              ways_3_metas_82_mru <= 1'b1;
            end
            if(_zz_1246) begin
              ways_3_metas_83_mru <= 1'b1;
            end
            if(_zz_1247) begin
              ways_3_metas_84_mru <= 1'b1;
            end
            if(_zz_1248) begin
              ways_3_metas_85_mru <= 1'b1;
            end
            if(_zz_1249) begin
              ways_3_metas_86_mru <= 1'b1;
            end
            if(_zz_1250) begin
              ways_3_metas_87_mru <= 1'b1;
            end
            if(_zz_1251) begin
              ways_3_metas_88_mru <= 1'b1;
            end
            if(_zz_1252) begin
              ways_3_metas_89_mru <= 1'b1;
            end
            if(_zz_1253) begin
              ways_3_metas_90_mru <= 1'b1;
            end
            if(_zz_1254) begin
              ways_3_metas_91_mru <= 1'b1;
            end
            if(_zz_1255) begin
              ways_3_metas_92_mru <= 1'b1;
            end
            if(_zz_1256) begin
              ways_3_metas_93_mru <= 1'b1;
            end
            if(_zz_1257) begin
              ways_3_metas_94_mru <= 1'b1;
            end
            if(_zz_1258) begin
              ways_3_metas_95_mru <= 1'b1;
            end
            if(_zz_1259) begin
              ways_3_metas_96_mru <= 1'b1;
            end
            if(_zz_1260) begin
              ways_3_metas_97_mru <= 1'b1;
            end
            if(_zz_1261) begin
              ways_3_metas_98_mru <= 1'b1;
            end
            if(_zz_1262) begin
              ways_3_metas_99_mru <= 1'b1;
            end
            if(_zz_1263) begin
              ways_3_metas_100_mru <= 1'b1;
            end
            if(_zz_1264) begin
              ways_3_metas_101_mru <= 1'b1;
            end
            if(_zz_1265) begin
              ways_3_metas_102_mru <= 1'b1;
            end
            if(_zz_1266) begin
              ways_3_metas_103_mru <= 1'b1;
            end
            if(_zz_1267) begin
              ways_3_metas_104_mru <= 1'b1;
            end
            if(_zz_1268) begin
              ways_3_metas_105_mru <= 1'b1;
            end
            if(_zz_1269) begin
              ways_3_metas_106_mru <= 1'b1;
            end
            if(_zz_1270) begin
              ways_3_metas_107_mru <= 1'b1;
            end
            if(_zz_1271) begin
              ways_3_metas_108_mru <= 1'b1;
            end
            if(_zz_1272) begin
              ways_3_metas_109_mru <= 1'b1;
            end
            if(_zz_1273) begin
              ways_3_metas_110_mru <= 1'b1;
            end
            if(_zz_1274) begin
              ways_3_metas_111_mru <= 1'b1;
            end
            if(_zz_1275) begin
              ways_3_metas_112_mru <= 1'b1;
            end
            if(_zz_1276) begin
              ways_3_metas_113_mru <= 1'b1;
            end
            if(_zz_1277) begin
              ways_3_metas_114_mru <= 1'b1;
            end
            if(_zz_1278) begin
              ways_3_metas_115_mru <= 1'b1;
            end
            if(_zz_1279) begin
              ways_3_metas_116_mru <= 1'b1;
            end
            if(_zz_1280) begin
              ways_3_metas_117_mru <= 1'b1;
            end
            if(_zz_1281) begin
              ways_3_metas_118_mru <= 1'b1;
            end
            if(_zz_1282) begin
              ways_3_metas_119_mru <= 1'b1;
            end
            if(_zz_1283) begin
              ways_3_metas_120_mru <= 1'b1;
            end
            if(_zz_1284) begin
              ways_3_metas_121_mru <= 1'b1;
            end
            if(_zz_1285) begin
              ways_3_metas_122_mru <= 1'b1;
            end
            if(_zz_1286) begin
              ways_3_metas_123_mru <= 1'b1;
            end
            if(_zz_1287) begin
              ways_3_metas_124_mru <= 1'b1;
            end
            if(_zz_1288) begin
              ways_3_metas_125_mru <= 1'b1;
            end
            if(_zz_1289) begin
              ways_3_metas_126_mru <= 1'b1;
            end
            if(_zz_1290) begin
              ways_3_metas_127_mru <= 1'b1;
            end
          end else begin
            if(when_ICache_l220_3) begin
              if(_zz_1292) begin
                ways_3_metas_0_vld <= 1'b1;
              end
              if(_zz_1293) begin
                ways_3_metas_1_vld <= 1'b1;
              end
              if(_zz_1294) begin
                ways_3_metas_2_vld <= 1'b1;
              end
              if(_zz_1295) begin
                ways_3_metas_3_vld <= 1'b1;
              end
              if(_zz_1296) begin
                ways_3_metas_4_vld <= 1'b1;
              end
              if(_zz_1297) begin
                ways_3_metas_5_vld <= 1'b1;
              end
              if(_zz_1298) begin
                ways_3_metas_6_vld <= 1'b1;
              end
              if(_zz_1299) begin
                ways_3_metas_7_vld <= 1'b1;
              end
              if(_zz_1300) begin
                ways_3_metas_8_vld <= 1'b1;
              end
              if(_zz_1301) begin
                ways_3_metas_9_vld <= 1'b1;
              end
              if(_zz_1302) begin
                ways_3_metas_10_vld <= 1'b1;
              end
              if(_zz_1303) begin
                ways_3_metas_11_vld <= 1'b1;
              end
              if(_zz_1304) begin
                ways_3_metas_12_vld <= 1'b1;
              end
              if(_zz_1305) begin
                ways_3_metas_13_vld <= 1'b1;
              end
              if(_zz_1306) begin
                ways_3_metas_14_vld <= 1'b1;
              end
              if(_zz_1307) begin
                ways_3_metas_15_vld <= 1'b1;
              end
              if(_zz_1308) begin
                ways_3_metas_16_vld <= 1'b1;
              end
              if(_zz_1309) begin
                ways_3_metas_17_vld <= 1'b1;
              end
              if(_zz_1310) begin
                ways_3_metas_18_vld <= 1'b1;
              end
              if(_zz_1311) begin
                ways_3_metas_19_vld <= 1'b1;
              end
              if(_zz_1312) begin
                ways_3_metas_20_vld <= 1'b1;
              end
              if(_zz_1313) begin
                ways_3_metas_21_vld <= 1'b1;
              end
              if(_zz_1314) begin
                ways_3_metas_22_vld <= 1'b1;
              end
              if(_zz_1315) begin
                ways_3_metas_23_vld <= 1'b1;
              end
              if(_zz_1316) begin
                ways_3_metas_24_vld <= 1'b1;
              end
              if(_zz_1317) begin
                ways_3_metas_25_vld <= 1'b1;
              end
              if(_zz_1318) begin
                ways_3_metas_26_vld <= 1'b1;
              end
              if(_zz_1319) begin
                ways_3_metas_27_vld <= 1'b1;
              end
              if(_zz_1320) begin
                ways_3_metas_28_vld <= 1'b1;
              end
              if(_zz_1321) begin
                ways_3_metas_29_vld <= 1'b1;
              end
              if(_zz_1322) begin
                ways_3_metas_30_vld <= 1'b1;
              end
              if(_zz_1323) begin
                ways_3_metas_31_vld <= 1'b1;
              end
              if(_zz_1324) begin
                ways_3_metas_32_vld <= 1'b1;
              end
              if(_zz_1325) begin
                ways_3_metas_33_vld <= 1'b1;
              end
              if(_zz_1326) begin
                ways_3_metas_34_vld <= 1'b1;
              end
              if(_zz_1327) begin
                ways_3_metas_35_vld <= 1'b1;
              end
              if(_zz_1328) begin
                ways_3_metas_36_vld <= 1'b1;
              end
              if(_zz_1329) begin
                ways_3_metas_37_vld <= 1'b1;
              end
              if(_zz_1330) begin
                ways_3_metas_38_vld <= 1'b1;
              end
              if(_zz_1331) begin
                ways_3_metas_39_vld <= 1'b1;
              end
              if(_zz_1332) begin
                ways_3_metas_40_vld <= 1'b1;
              end
              if(_zz_1333) begin
                ways_3_metas_41_vld <= 1'b1;
              end
              if(_zz_1334) begin
                ways_3_metas_42_vld <= 1'b1;
              end
              if(_zz_1335) begin
                ways_3_metas_43_vld <= 1'b1;
              end
              if(_zz_1336) begin
                ways_3_metas_44_vld <= 1'b1;
              end
              if(_zz_1337) begin
                ways_3_metas_45_vld <= 1'b1;
              end
              if(_zz_1338) begin
                ways_3_metas_46_vld <= 1'b1;
              end
              if(_zz_1339) begin
                ways_3_metas_47_vld <= 1'b1;
              end
              if(_zz_1340) begin
                ways_3_metas_48_vld <= 1'b1;
              end
              if(_zz_1341) begin
                ways_3_metas_49_vld <= 1'b1;
              end
              if(_zz_1342) begin
                ways_3_metas_50_vld <= 1'b1;
              end
              if(_zz_1343) begin
                ways_3_metas_51_vld <= 1'b1;
              end
              if(_zz_1344) begin
                ways_3_metas_52_vld <= 1'b1;
              end
              if(_zz_1345) begin
                ways_3_metas_53_vld <= 1'b1;
              end
              if(_zz_1346) begin
                ways_3_metas_54_vld <= 1'b1;
              end
              if(_zz_1347) begin
                ways_3_metas_55_vld <= 1'b1;
              end
              if(_zz_1348) begin
                ways_3_metas_56_vld <= 1'b1;
              end
              if(_zz_1349) begin
                ways_3_metas_57_vld <= 1'b1;
              end
              if(_zz_1350) begin
                ways_3_metas_58_vld <= 1'b1;
              end
              if(_zz_1351) begin
                ways_3_metas_59_vld <= 1'b1;
              end
              if(_zz_1352) begin
                ways_3_metas_60_vld <= 1'b1;
              end
              if(_zz_1353) begin
                ways_3_metas_61_vld <= 1'b1;
              end
              if(_zz_1354) begin
                ways_3_metas_62_vld <= 1'b1;
              end
              if(_zz_1355) begin
                ways_3_metas_63_vld <= 1'b1;
              end
              if(_zz_1356) begin
                ways_3_metas_64_vld <= 1'b1;
              end
              if(_zz_1357) begin
                ways_3_metas_65_vld <= 1'b1;
              end
              if(_zz_1358) begin
                ways_3_metas_66_vld <= 1'b1;
              end
              if(_zz_1359) begin
                ways_3_metas_67_vld <= 1'b1;
              end
              if(_zz_1360) begin
                ways_3_metas_68_vld <= 1'b1;
              end
              if(_zz_1361) begin
                ways_3_metas_69_vld <= 1'b1;
              end
              if(_zz_1362) begin
                ways_3_metas_70_vld <= 1'b1;
              end
              if(_zz_1363) begin
                ways_3_metas_71_vld <= 1'b1;
              end
              if(_zz_1364) begin
                ways_3_metas_72_vld <= 1'b1;
              end
              if(_zz_1365) begin
                ways_3_metas_73_vld <= 1'b1;
              end
              if(_zz_1366) begin
                ways_3_metas_74_vld <= 1'b1;
              end
              if(_zz_1367) begin
                ways_3_metas_75_vld <= 1'b1;
              end
              if(_zz_1368) begin
                ways_3_metas_76_vld <= 1'b1;
              end
              if(_zz_1369) begin
                ways_3_metas_77_vld <= 1'b1;
              end
              if(_zz_1370) begin
                ways_3_metas_78_vld <= 1'b1;
              end
              if(_zz_1371) begin
                ways_3_metas_79_vld <= 1'b1;
              end
              if(_zz_1372) begin
                ways_3_metas_80_vld <= 1'b1;
              end
              if(_zz_1373) begin
                ways_3_metas_81_vld <= 1'b1;
              end
              if(_zz_1374) begin
                ways_3_metas_82_vld <= 1'b1;
              end
              if(_zz_1375) begin
                ways_3_metas_83_vld <= 1'b1;
              end
              if(_zz_1376) begin
                ways_3_metas_84_vld <= 1'b1;
              end
              if(_zz_1377) begin
                ways_3_metas_85_vld <= 1'b1;
              end
              if(_zz_1378) begin
                ways_3_metas_86_vld <= 1'b1;
              end
              if(_zz_1379) begin
                ways_3_metas_87_vld <= 1'b1;
              end
              if(_zz_1380) begin
                ways_3_metas_88_vld <= 1'b1;
              end
              if(_zz_1381) begin
                ways_3_metas_89_vld <= 1'b1;
              end
              if(_zz_1382) begin
                ways_3_metas_90_vld <= 1'b1;
              end
              if(_zz_1383) begin
                ways_3_metas_91_vld <= 1'b1;
              end
              if(_zz_1384) begin
                ways_3_metas_92_vld <= 1'b1;
              end
              if(_zz_1385) begin
                ways_3_metas_93_vld <= 1'b1;
              end
              if(_zz_1386) begin
                ways_3_metas_94_vld <= 1'b1;
              end
              if(_zz_1387) begin
                ways_3_metas_95_vld <= 1'b1;
              end
              if(_zz_1388) begin
                ways_3_metas_96_vld <= 1'b1;
              end
              if(_zz_1389) begin
                ways_3_metas_97_vld <= 1'b1;
              end
              if(_zz_1390) begin
                ways_3_metas_98_vld <= 1'b1;
              end
              if(_zz_1391) begin
                ways_3_metas_99_vld <= 1'b1;
              end
              if(_zz_1392) begin
                ways_3_metas_100_vld <= 1'b1;
              end
              if(_zz_1393) begin
                ways_3_metas_101_vld <= 1'b1;
              end
              if(_zz_1394) begin
                ways_3_metas_102_vld <= 1'b1;
              end
              if(_zz_1395) begin
                ways_3_metas_103_vld <= 1'b1;
              end
              if(_zz_1396) begin
                ways_3_metas_104_vld <= 1'b1;
              end
              if(_zz_1397) begin
                ways_3_metas_105_vld <= 1'b1;
              end
              if(_zz_1398) begin
                ways_3_metas_106_vld <= 1'b1;
              end
              if(_zz_1399) begin
                ways_3_metas_107_vld <= 1'b1;
              end
              if(_zz_1400) begin
                ways_3_metas_108_vld <= 1'b1;
              end
              if(_zz_1401) begin
                ways_3_metas_109_vld <= 1'b1;
              end
              if(_zz_1402) begin
                ways_3_metas_110_vld <= 1'b1;
              end
              if(_zz_1403) begin
                ways_3_metas_111_vld <= 1'b1;
              end
              if(_zz_1404) begin
                ways_3_metas_112_vld <= 1'b1;
              end
              if(_zz_1405) begin
                ways_3_metas_113_vld <= 1'b1;
              end
              if(_zz_1406) begin
                ways_3_metas_114_vld <= 1'b1;
              end
              if(_zz_1407) begin
                ways_3_metas_115_vld <= 1'b1;
              end
              if(_zz_1408) begin
                ways_3_metas_116_vld <= 1'b1;
              end
              if(_zz_1409) begin
                ways_3_metas_117_vld <= 1'b1;
              end
              if(_zz_1410) begin
                ways_3_metas_118_vld <= 1'b1;
              end
              if(_zz_1411) begin
                ways_3_metas_119_vld <= 1'b1;
              end
              if(_zz_1412) begin
                ways_3_metas_120_vld <= 1'b1;
              end
              if(_zz_1413) begin
                ways_3_metas_121_vld <= 1'b1;
              end
              if(_zz_1414) begin
                ways_3_metas_122_vld <= 1'b1;
              end
              if(_zz_1415) begin
                ways_3_metas_123_vld <= 1'b1;
              end
              if(_zz_1416) begin
                ways_3_metas_124_vld <= 1'b1;
              end
              if(_zz_1417) begin
                ways_3_metas_125_vld <= 1'b1;
              end
              if(_zz_1418) begin
                ways_3_metas_126_vld <= 1'b1;
              end
              if(_zz_1419) begin
                ways_3_metas_127_vld <= 1'b1;
              end
            end
          end
        end
      end
      if(when_ICache_l225_3) begin
        if(_zz_1292) begin
          ways_3_metas_0_tag <= cpu_tag_d1;
        end
        if(_zz_1293) begin
          ways_3_metas_1_tag <= cpu_tag_d1;
        end
        if(_zz_1294) begin
          ways_3_metas_2_tag <= cpu_tag_d1;
        end
        if(_zz_1295) begin
          ways_3_metas_3_tag <= cpu_tag_d1;
        end
        if(_zz_1296) begin
          ways_3_metas_4_tag <= cpu_tag_d1;
        end
        if(_zz_1297) begin
          ways_3_metas_5_tag <= cpu_tag_d1;
        end
        if(_zz_1298) begin
          ways_3_metas_6_tag <= cpu_tag_d1;
        end
        if(_zz_1299) begin
          ways_3_metas_7_tag <= cpu_tag_d1;
        end
        if(_zz_1300) begin
          ways_3_metas_8_tag <= cpu_tag_d1;
        end
        if(_zz_1301) begin
          ways_3_metas_9_tag <= cpu_tag_d1;
        end
        if(_zz_1302) begin
          ways_3_metas_10_tag <= cpu_tag_d1;
        end
        if(_zz_1303) begin
          ways_3_metas_11_tag <= cpu_tag_d1;
        end
        if(_zz_1304) begin
          ways_3_metas_12_tag <= cpu_tag_d1;
        end
        if(_zz_1305) begin
          ways_3_metas_13_tag <= cpu_tag_d1;
        end
        if(_zz_1306) begin
          ways_3_metas_14_tag <= cpu_tag_d1;
        end
        if(_zz_1307) begin
          ways_3_metas_15_tag <= cpu_tag_d1;
        end
        if(_zz_1308) begin
          ways_3_metas_16_tag <= cpu_tag_d1;
        end
        if(_zz_1309) begin
          ways_3_metas_17_tag <= cpu_tag_d1;
        end
        if(_zz_1310) begin
          ways_3_metas_18_tag <= cpu_tag_d1;
        end
        if(_zz_1311) begin
          ways_3_metas_19_tag <= cpu_tag_d1;
        end
        if(_zz_1312) begin
          ways_3_metas_20_tag <= cpu_tag_d1;
        end
        if(_zz_1313) begin
          ways_3_metas_21_tag <= cpu_tag_d1;
        end
        if(_zz_1314) begin
          ways_3_metas_22_tag <= cpu_tag_d1;
        end
        if(_zz_1315) begin
          ways_3_metas_23_tag <= cpu_tag_d1;
        end
        if(_zz_1316) begin
          ways_3_metas_24_tag <= cpu_tag_d1;
        end
        if(_zz_1317) begin
          ways_3_metas_25_tag <= cpu_tag_d1;
        end
        if(_zz_1318) begin
          ways_3_metas_26_tag <= cpu_tag_d1;
        end
        if(_zz_1319) begin
          ways_3_metas_27_tag <= cpu_tag_d1;
        end
        if(_zz_1320) begin
          ways_3_metas_28_tag <= cpu_tag_d1;
        end
        if(_zz_1321) begin
          ways_3_metas_29_tag <= cpu_tag_d1;
        end
        if(_zz_1322) begin
          ways_3_metas_30_tag <= cpu_tag_d1;
        end
        if(_zz_1323) begin
          ways_3_metas_31_tag <= cpu_tag_d1;
        end
        if(_zz_1324) begin
          ways_3_metas_32_tag <= cpu_tag_d1;
        end
        if(_zz_1325) begin
          ways_3_metas_33_tag <= cpu_tag_d1;
        end
        if(_zz_1326) begin
          ways_3_metas_34_tag <= cpu_tag_d1;
        end
        if(_zz_1327) begin
          ways_3_metas_35_tag <= cpu_tag_d1;
        end
        if(_zz_1328) begin
          ways_3_metas_36_tag <= cpu_tag_d1;
        end
        if(_zz_1329) begin
          ways_3_metas_37_tag <= cpu_tag_d1;
        end
        if(_zz_1330) begin
          ways_3_metas_38_tag <= cpu_tag_d1;
        end
        if(_zz_1331) begin
          ways_3_metas_39_tag <= cpu_tag_d1;
        end
        if(_zz_1332) begin
          ways_3_metas_40_tag <= cpu_tag_d1;
        end
        if(_zz_1333) begin
          ways_3_metas_41_tag <= cpu_tag_d1;
        end
        if(_zz_1334) begin
          ways_3_metas_42_tag <= cpu_tag_d1;
        end
        if(_zz_1335) begin
          ways_3_metas_43_tag <= cpu_tag_d1;
        end
        if(_zz_1336) begin
          ways_3_metas_44_tag <= cpu_tag_d1;
        end
        if(_zz_1337) begin
          ways_3_metas_45_tag <= cpu_tag_d1;
        end
        if(_zz_1338) begin
          ways_3_metas_46_tag <= cpu_tag_d1;
        end
        if(_zz_1339) begin
          ways_3_metas_47_tag <= cpu_tag_d1;
        end
        if(_zz_1340) begin
          ways_3_metas_48_tag <= cpu_tag_d1;
        end
        if(_zz_1341) begin
          ways_3_metas_49_tag <= cpu_tag_d1;
        end
        if(_zz_1342) begin
          ways_3_metas_50_tag <= cpu_tag_d1;
        end
        if(_zz_1343) begin
          ways_3_metas_51_tag <= cpu_tag_d1;
        end
        if(_zz_1344) begin
          ways_3_metas_52_tag <= cpu_tag_d1;
        end
        if(_zz_1345) begin
          ways_3_metas_53_tag <= cpu_tag_d1;
        end
        if(_zz_1346) begin
          ways_3_metas_54_tag <= cpu_tag_d1;
        end
        if(_zz_1347) begin
          ways_3_metas_55_tag <= cpu_tag_d1;
        end
        if(_zz_1348) begin
          ways_3_metas_56_tag <= cpu_tag_d1;
        end
        if(_zz_1349) begin
          ways_3_metas_57_tag <= cpu_tag_d1;
        end
        if(_zz_1350) begin
          ways_3_metas_58_tag <= cpu_tag_d1;
        end
        if(_zz_1351) begin
          ways_3_metas_59_tag <= cpu_tag_d1;
        end
        if(_zz_1352) begin
          ways_3_metas_60_tag <= cpu_tag_d1;
        end
        if(_zz_1353) begin
          ways_3_metas_61_tag <= cpu_tag_d1;
        end
        if(_zz_1354) begin
          ways_3_metas_62_tag <= cpu_tag_d1;
        end
        if(_zz_1355) begin
          ways_3_metas_63_tag <= cpu_tag_d1;
        end
        if(_zz_1356) begin
          ways_3_metas_64_tag <= cpu_tag_d1;
        end
        if(_zz_1357) begin
          ways_3_metas_65_tag <= cpu_tag_d1;
        end
        if(_zz_1358) begin
          ways_3_metas_66_tag <= cpu_tag_d1;
        end
        if(_zz_1359) begin
          ways_3_metas_67_tag <= cpu_tag_d1;
        end
        if(_zz_1360) begin
          ways_3_metas_68_tag <= cpu_tag_d1;
        end
        if(_zz_1361) begin
          ways_3_metas_69_tag <= cpu_tag_d1;
        end
        if(_zz_1362) begin
          ways_3_metas_70_tag <= cpu_tag_d1;
        end
        if(_zz_1363) begin
          ways_3_metas_71_tag <= cpu_tag_d1;
        end
        if(_zz_1364) begin
          ways_3_metas_72_tag <= cpu_tag_d1;
        end
        if(_zz_1365) begin
          ways_3_metas_73_tag <= cpu_tag_d1;
        end
        if(_zz_1366) begin
          ways_3_metas_74_tag <= cpu_tag_d1;
        end
        if(_zz_1367) begin
          ways_3_metas_75_tag <= cpu_tag_d1;
        end
        if(_zz_1368) begin
          ways_3_metas_76_tag <= cpu_tag_d1;
        end
        if(_zz_1369) begin
          ways_3_metas_77_tag <= cpu_tag_d1;
        end
        if(_zz_1370) begin
          ways_3_metas_78_tag <= cpu_tag_d1;
        end
        if(_zz_1371) begin
          ways_3_metas_79_tag <= cpu_tag_d1;
        end
        if(_zz_1372) begin
          ways_3_metas_80_tag <= cpu_tag_d1;
        end
        if(_zz_1373) begin
          ways_3_metas_81_tag <= cpu_tag_d1;
        end
        if(_zz_1374) begin
          ways_3_metas_82_tag <= cpu_tag_d1;
        end
        if(_zz_1375) begin
          ways_3_metas_83_tag <= cpu_tag_d1;
        end
        if(_zz_1376) begin
          ways_3_metas_84_tag <= cpu_tag_d1;
        end
        if(_zz_1377) begin
          ways_3_metas_85_tag <= cpu_tag_d1;
        end
        if(_zz_1378) begin
          ways_3_metas_86_tag <= cpu_tag_d1;
        end
        if(_zz_1379) begin
          ways_3_metas_87_tag <= cpu_tag_d1;
        end
        if(_zz_1380) begin
          ways_3_metas_88_tag <= cpu_tag_d1;
        end
        if(_zz_1381) begin
          ways_3_metas_89_tag <= cpu_tag_d1;
        end
        if(_zz_1382) begin
          ways_3_metas_90_tag <= cpu_tag_d1;
        end
        if(_zz_1383) begin
          ways_3_metas_91_tag <= cpu_tag_d1;
        end
        if(_zz_1384) begin
          ways_3_metas_92_tag <= cpu_tag_d1;
        end
        if(_zz_1385) begin
          ways_3_metas_93_tag <= cpu_tag_d1;
        end
        if(_zz_1386) begin
          ways_3_metas_94_tag <= cpu_tag_d1;
        end
        if(_zz_1387) begin
          ways_3_metas_95_tag <= cpu_tag_d1;
        end
        if(_zz_1388) begin
          ways_3_metas_96_tag <= cpu_tag_d1;
        end
        if(_zz_1389) begin
          ways_3_metas_97_tag <= cpu_tag_d1;
        end
        if(_zz_1390) begin
          ways_3_metas_98_tag <= cpu_tag_d1;
        end
        if(_zz_1391) begin
          ways_3_metas_99_tag <= cpu_tag_d1;
        end
        if(_zz_1392) begin
          ways_3_metas_100_tag <= cpu_tag_d1;
        end
        if(_zz_1393) begin
          ways_3_metas_101_tag <= cpu_tag_d1;
        end
        if(_zz_1394) begin
          ways_3_metas_102_tag <= cpu_tag_d1;
        end
        if(_zz_1395) begin
          ways_3_metas_103_tag <= cpu_tag_d1;
        end
        if(_zz_1396) begin
          ways_3_metas_104_tag <= cpu_tag_d1;
        end
        if(_zz_1397) begin
          ways_3_metas_105_tag <= cpu_tag_d1;
        end
        if(_zz_1398) begin
          ways_3_metas_106_tag <= cpu_tag_d1;
        end
        if(_zz_1399) begin
          ways_3_metas_107_tag <= cpu_tag_d1;
        end
        if(_zz_1400) begin
          ways_3_metas_108_tag <= cpu_tag_d1;
        end
        if(_zz_1401) begin
          ways_3_metas_109_tag <= cpu_tag_d1;
        end
        if(_zz_1402) begin
          ways_3_metas_110_tag <= cpu_tag_d1;
        end
        if(_zz_1403) begin
          ways_3_metas_111_tag <= cpu_tag_d1;
        end
        if(_zz_1404) begin
          ways_3_metas_112_tag <= cpu_tag_d1;
        end
        if(_zz_1405) begin
          ways_3_metas_113_tag <= cpu_tag_d1;
        end
        if(_zz_1406) begin
          ways_3_metas_114_tag <= cpu_tag_d1;
        end
        if(_zz_1407) begin
          ways_3_metas_115_tag <= cpu_tag_d1;
        end
        if(_zz_1408) begin
          ways_3_metas_116_tag <= cpu_tag_d1;
        end
        if(_zz_1409) begin
          ways_3_metas_117_tag <= cpu_tag_d1;
        end
        if(_zz_1410) begin
          ways_3_metas_118_tag <= cpu_tag_d1;
        end
        if(_zz_1411) begin
          ways_3_metas_119_tag <= cpu_tag_d1;
        end
        if(_zz_1412) begin
          ways_3_metas_120_tag <= cpu_tag_d1;
        end
        if(_zz_1413) begin
          ways_3_metas_121_tag <= cpu_tag_d1;
        end
        if(_zz_1414) begin
          ways_3_metas_122_tag <= cpu_tag_d1;
        end
        if(_zz_1415) begin
          ways_3_metas_123_tag <= cpu_tag_d1;
        end
        if(_zz_1416) begin
          ways_3_metas_124_tag <= cpu_tag_d1;
        end
        if(_zz_1417) begin
          ways_3_metas_125_tag <= cpu_tag_d1;
        end
        if(_zz_1418) begin
          ways_3_metas_126_tag <= cpu_tag_d1;
        end
        if(_zz_1419) begin
          ways_3_metas_127_tag <= cpu_tag_d1;
        end
      end
      if(when_ICache_l230_3) begin
        cpu_cmd_ready_1 <= 1'b0;
      end else begin
        if(when_ICache_l233_3) begin
          cpu_cmd_ready_1 <= 1'b1;
        end
      end
    end
  end

  always @(posedge clk) begin
    hit_id_d1 <= hit_id;
    is_hit_d1 <= is_hit;
    if(is_miss) begin
      evict_id_miss <= evict_id;
    end
    next_level_done <= (next_level_rsp_valid && (next_level_data_cnt_value == 3'b111));
  end


endmodule

module Timer (
  input               cen,
  input               wen,
  input      [63:0]   addr,
  input      [63:0]   wdata,
  output reg [63:0]   rdata,
  output              timer_int,
  input               clk,
  input               reset
);

  wire       [63:0]   _zz_mtime;
  reg        [63:0]   mtime;
  reg        [63:0]   mtimecmp;
  wire                when_ExcepPlugin_l277;
  wire                when_ExcepPlugin_l290;
  wire                when_ExcepPlugin_l292;

  assign _zz_mtime = (mtime + 64'h0000000000000001);
  assign when_ExcepPlugin_l277 = (wen && cen);
  assign when_ExcepPlugin_l290 = (addr == 64'h000000000200bff8);
  always @(*) begin
    if(when_ExcepPlugin_l290) begin
      rdata = mtime;
    end else begin
      if(when_ExcepPlugin_l292) begin
        rdata = mtimecmp;
      end else begin
        rdata = 64'h0;
      end
    end
  end

  assign when_ExcepPlugin_l292 = (addr == 64'h0000000002004000);
  assign timer_int = (mtimecmp <= mtime);
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      mtime <= 64'h0;
      mtimecmp <= 64'hffffffffffffffff;
    end else begin
      if(when_ExcepPlugin_l277) begin
        case(addr)
          64'h000000000200bff8 : begin
            mtime <= wdata;
          end
          64'h0000000002004000 : begin
            mtimecmp <= wdata;
          end
          default : begin
          end
        endcase
      end else begin
        mtime <= _zz_mtime;
      end
    end
  end


endmodule

module Clint (
  input      [63:0]   pc,
  input      [63:0]   pc_next,
  input               pc_next_valid,
  input               instruction_valid,
  output reg          csr_ports_mepc_wen,
  output reg [63:0]   csr_ports_mepc_wdata,
  output reg          csr_ports_mcause_wen,
  output reg [63:0]   csr_ports_mcause_wdata,
  output reg          csr_ports_mstatus_wen,
  output reg [63:0]   csr_ports_mstatus_wdata,
  input      [63:0]   csr_ports_mtvec,
  input      [63:0]   csr_ports_mepc,
  input      [63:0]   csr_ports_mstatus,
  input               csr_ports_global_int_en,
  input               csr_ports_mtime_int_en,
  input               csr_ports_mtime_int_pend,
  input               timer_int,
  output reg          int_en,
  output reg [63:0]   int_pc,
  output              int_hold,
  input               ecall,
  input               ebreak,
  input               mret,
  input               clk,
  input               reset
);
  localparam IntTypeEnum_IDLE = 2'd0;
  localparam IntTypeEnum_EXPT = 2'd1;
  localparam IntTypeEnum_TIME_1 = 2'd2;
  localparam IntTypeEnum_MRET = 2'd3;

  reg        [1:0]    int_state;
  reg        [63:0]   pc_next_d1;
  reg        [63:0]   mepc_wdata;
  reg        [63:0]   mcause_wdata;
  wire                when_ExcepPlugin_l180;
  wire                when_ExcepPlugin_l182;
  wire                when_ExcepPlugin_l191;
  wire                when_ExcepPlugin_l208;
  wire                when_ExcepPlugin_l216;

  assign when_ExcepPlugin_l180 = (ecall || ebreak);
  always @(*) begin
    if(when_ExcepPlugin_l180) begin
      int_state = IntTypeEnum_EXPT;
    end else begin
      if(when_ExcepPlugin_l182) begin
        int_state = IntTypeEnum_TIME_1;
      end else begin
        if(mret) begin
          int_state = IntTypeEnum_MRET;
        end else begin
          int_state = IntTypeEnum_IDLE;
        end
      end
    end
  end

  assign when_ExcepPlugin_l182 = ((csr_ports_global_int_en && csr_ports_mtime_int_en) && timer_int);
  assign when_ExcepPlugin_l191 = (int_state == IntTypeEnum_TIME_1);
  always @(*) begin
    if(when_ExcepPlugin_l191) begin
      if(instruction_valid) begin
        mepc_wdata = pc_next;
      end else begin
        mepc_wdata = pc_next_d1;
      end
    end else begin
      if(instruction_valid) begin
        mepc_wdata = pc;
      end else begin
        mepc_wdata = pc_next_d1;
      end
    end
  end

  assign when_ExcepPlugin_l208 = (int_state == IntTypeEnum_EXPT);
  always @(*) begin
    if(when_ExcepPlugin_l208) begin
      if(ecall) begin
        mcause_wdata = 64'h000000000000000b;
      end else begin
        if(ebreak) begin
          mcause_wdata = 64'h0000000000000003;
        end else begin
          mcause_wdata = 64'h000000000000000a;
        end
      end
    end else begin
      if(when_ExcepPlugin_l216) begin
        mcause_wdata = 64'h8000000000000007;
      end else begin
        mcause_wdata = 64'h0;
      end
    end
  end

  assign when_ExcepPlugin_l216 = (int_state == IntTypeEnum_TIME_1);
  always @(*) begin
    if((int_state == IntTypeEnum_EXPT) || (int_state == IntTypeEnum_TIME_1)) begin
        int_en = 1'b1;
    end else if((int_state == IntTypeEnum_MRET)) begin
        int_en = 1'b1;
    end else begin
        int_en = 1'b0;
    end
  end

  always @(*) begin
    if((int_state == IntTypeEnum_EXPT) || (int_state == IntTypeEnum_TIME_1)) begin
        int_pc = csr_ports_mtvec;
    end else if((int_state == IntTypeEnum_MRET)) begin
        int_pc = csr_ports_mepc;
    end else begin
        int_pc = 64'h0;
    end
  end

  always @(*) begin
    if((int_state == IntTypeEnum_EXPT) || (int_state == IntTypeEnum_TIME_1)) begin
        csr_ports_mepc_wen = 1'b1;
    end else if((int_state == IntTypeEnum_MRET)) begin
        csr_ports_mepc_wen = 1'b0;
    end else begin
        csr_ports_mepc_wen = 1'b0;
    end
  end

  always @(*) begin
    if((int_state == IntTypeEnum_EXPT) || (int_state == IntTypeEnum_TIME_1)) begin
        csr_ports_mcause_wen = 1'b1;
    end else if((int_state == IntTypeEnum_MRET)) begin
        csr_ports_mcause_wen = 1'b0;
    end else begin
        csr_ports_mcause_wen = 1'b0;
    end
  end

  always @(*) begin
    if((int_state == IntTypeEnum_EXPT) || (int_state == IntTypeEnum_TIME_1)) begin
        csr_ports_mstatus_wen = 1'b1;
    end else if((int_state == IntTypeEnum_MRET)) begin
        csr_ports_mstatus_wen = 1'b1;
    end else begin
        csr_ports_mstatus_wen = 1'b0;
    end
  end

  always @(*) begin
    if((int_state == IntTypeEnum_EXPT) || (int_state == IntTypeEnum_TIME_1)) begin
        csr_ports_mepc_wdata = mepc_wdata;
    end else if((int_state == IntTypeEnum_MRET)) begin
        csr_ports_mepc_wdata = 64'h0;
    end else begin
        csr_ports_mepc_wdata = 64'h0;
    end
  end

  always @(*) begin
    if((int_state == IntTypeEnum_EXPT) || (int_state == IntTypeEnum_TIME_1)) begin
        csr_ports_mcause_wdata = mcause_wdata;
    end else if((int_state == IntTypeEnum_MRET)) begin
        csr_ports_mcause_wdata = 64'h0;
    end else begin
        csr_ports_mcause_wdata = 64'h0;
    end
  end

  always @(*) begin
    if((int_state == IntTypeEnum_EXPT) || (int_state == IntTypeEnum_TIME_1)) begin
        csr_ports_mstatus_wdata = {{{{csr_ports_mstatus[63 : 8],csr_ports_mstatus[3]},csr_ports_mstatus[6 : 4]},1'b0},csr_ports_mstatus[2 : 0]};
    end else if((int_state == IntTypeEnum_MRET)) begin
        csr_ports_mstatus_wdata = {{{{csr_ports_mstatus[63 : 8],1'b1},csr_ports_mstatus[6 : 4]},csr_ports_mstatus[7]},csr_ports_mstatus[2 : 0]};
    end else begin
        csr_ports_mstatus_wdata = 64'h0;
    end
  end

  assign int_hold = 1'b0;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      pc_next_d1 <= 64'h0;
    end else begin
      if(pc_next_valid) begin
        pc_next_d1 <= pc_next;
      end
    end
  end


endmodule

module CsrRegfile (
  input      [11:0]   cpu_ports_waddr,
  input               cpu_ports_wen,
  input      [63:0]   cpu_ports_wdata,
  input      [11:0]   cpu_ports_raddr,
  output reg [63:0]   cpu_ports_rdata,
  input               clint_ports_mepc_wen,
  input      [63:0]   clint_ports_mepc_wdata,
  input               clint_ports_mcause_wen,
  input      [63:0]   clint_ports_mcause_wdata,
  input               clint_ports_mstatus_wen,
  input      [63:0]   clint_ports_mstatus_wdata,
  output     [63:0]   clint_ports_mtvec,
  output     [63:0]   clint_ports_mepc,
  output     [63:0]   clint_ports_mstatus,
  output              clint_ports_global_int_en,
  output              clint_ports_mtime_int_en,
  output              clint_ports_mtime_int_pend,
  input               timer_int,
  input               clk,
  input               reset
);

  wire       [63:0]   _zz_mcycle;
  reg        [63:0]   mstatus;
  reg        [63:0]   mie;
  reg        [63:0]   mtvec;
  reg        [63:0]   mepc;
  reg        [63:0]   mcause;
  reg        [63:0]   mtval;
  reg        [63:0]   mip;
  reg        [63:0]   mcycle;
  reg        [63:0]   mhartid;
  reg        [63:0]   mscratch;
  wire                when_ExcepPlugin_l106;

  assign _zz_mcycle = (mcycle + 64'h0000000000000001);
  assign when_ExcepPlugin_l106 = (cpu_ports_wen && (cpu_ports_raddr == cpu_ports_waddr));
  always @(*) begin
    if(when_ExcepPlugin_l106) begin
      cpu_ports_rdata = cpu_ports_wdata;
    end else begin
      case(cpu_ports_raddr)
        12'h300 : begin
          cpu_ports_rdata = mstatus;
        end
        12'h304 : begin
          cpu_ports_rdata = mie;
        end
        12'h305 : begin
          cpu_ports_rdata = mtvec;
        end
        12'h341 : begin
          cpu_ports_rdata = mepc;
        end
        12'h342 : begin
          cpu_ports_rdata = mcause;
        end
        12'h343 : begin
          cpu_ports_rdata = mtval;
        end
        12'h344 : begin
          cpu_ports_rdata = mip;
        end
        12'hb00 : begin
          cpu_ports_rdata = mcycle;
        end
        12'hf14 : begin
          cpu_ports_rdata = mhartid;
        end
        default : begin
          cpu_ports_rdata = 64'h0;
        end
      endcase
    end
  end

  assign clint_ports_mtvec = mtvec;
  assign clint_ports_mepc = mepc;
  assign clint_ports_mstatus = mstatus;
  assign clint_ports_global_int_en = mstatus[3];
  assign clint_ports_mtime_int_en = mie[7];
  assign clint_ports_mtime_int_pend = mip[7];
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      mstatus <= {51'h0,13'h1880};
      mie <= 64'h0;
      mtvec <= 64'h0;
      mepc <= 64'h0;
      mcause <= 64'h0;
      mtval <= 64'h0;
      mip <= 64'h0;
      mcycle <= 64'h0;
      mhartid <= 64'h0;
      mscratch <= 64'h0;
    end else begin
      mcycle <= _zz_mcycle;
      mip <= {{{{52'h0,1'b0},3'b000},timer_int},7'h0};
      if(cpu_ports_wen) begin
        case(cpu_ports_waddr)
          12'h300 : begin
            mstatus <= {{{{{{{((cpu_ports_wdata[16 : 15] == 2'b11) || (cpu_ports_wdata[14 : 13] == 2'b11)),50'h0},2'b11},3'b000},cpu_ports_wdata[7]},3'b000},cpu_ports_wdata[3]},3'b000};
          end
          12'h304 : begin
            mie <= {{{{{{52'h0,cpu_ports_wdata[11]},3'b000},cpu_ports_wdata[7]},3'b000},cpu_ports_wdata[3]},3'b000};
          end
          12'h305 : begin
            mtvec <= cpu_ports_wdata;
          end
          12'h341 : begin
            mepc <= cpu_ports_wdata;
          end
          12'h342 : begin
            mcause <= cpu_ports_wdata;
          end
          12'h343 : begin
            mtval <= cpu_ports_wdata;
          end
          12'hf14 : begin
            mhartid <= cpu_ports_wdata;
          end
          12'h340 : begin
            mscratch <= cpu_ports_wdata;
          end
          default : begin
          end
        endcase
      end else begin
        if(clint_ports_mepc_wen) begin
          mepc <= clint_ports_mepc_wdata;
        end
        if(clint_ports_mcause_wen) begin
          mcause <= clint_ports_mcause_wdata;
        end
        if(clint_ports_mstatus_wen) begin
          mstatus <= clint_ports_mstatus_wdata;
        end
        mtvec <= {clint_ports_mtvec[63 : 2],2'b00};
      end
    end
  end


endmodule

module RegFileModule (
  output     [63:0]   read_ports_rs1_value,
  output     [63:0]   read_ports_rs2_value,
  input      [4:0]    read_ports_rs1_addr,
  input      [4:0]    read_ports_rs2_addr,
  input               read_ports_rs1_req,
  input               read_ports_rs2_req,
  input      [63:0]   write_ports_rd_value,
  input      [4:0]    write_ports_rd_addr,
  input               write_ports_rd_wen,
  input               clk,
  input               reset
);

  reg        [63:0]   _zz_read_value_1;
  reg        [63:0]   _zz_read_value_2;
  reg        [63:0]   reg_file_0;
  reg        [63:0]   reg_file_1;
  reg        [63:0]   reg_file_2;
  reg        [63:0]   reg_file_3;
  reg        [63:0]   reg_file_4;
  reg        [63:0]   reg_file_5;
  reg        [63:0]   reg_file_6;
  reg        [63:0]   reg_file_7;
  reg        [63:0]   reg_file_8;
  reg        [63:0]   reg_file_9;
  reg        [63:0]   reg_file_10;
  reg        [63:0]   reg_file_11;
  reg        [63:0]   reg_file_12;
  reg        [63:0]   reg_file_13;
  reg        [63:0]   reg_file_14;
  reg        [63:0]   reg_file_15;
  reg        [63:0]   reg_file_16;
  reg        [63:0]   reg_file_17;
  reg        [63:0]   reg_file_18;
  reg        [63:0]   reg_file_19;
  reg        [63:0]   reg_file_20;
  reg        [63:0]   reg_file_21;
  reg        [63:0]   reg_file_22;
  reg        [63:0]   reg_file_23;
  reg        [63:0]   reg_file_24;
  reg        [63:0]   reg_file_25;
  reg        [63:0]   reg_file_26;
  reg        [63:0]   reg_file_27;
  reg        [63:0]   reg_file_28;
  reg        [63:0]   reg_file_29;
  reg        [63:0]   reg_file_30;
  reg        [63:0]   reg_file_31;
  wire       [63:0]   read_value_1;
  wire       [63:0]   read_value_2;
  wire                when_DecodePlugin_l61;
  wire       [31:0]   _zz_1;

  always @(*) begin
    case(read_ports_rs1_addr)
      5'b00000 : _zz_read_value_1 = reg_file_0;
      5'b00001 : _zz_read_value_1 = reg_file_1;
      5'b00010 : _zz_read_value_1 = reg_file_2;
      5'b00011 : _zz_read_value_1 = reg_file_3;
      5'b00100 : _zz_read_value_1 = reg_file_4;
      5'b00101 : _zz_read_value_1 = reg_file_5;
      5'b00110 : _zz_read_value_1 = reg_file_6;
      5'b00111 : _zz_read_value_1 = reg_file_7;
      5'b01000 : _zz_read_value_1 = reg_file_8;
      5'b01001 : _zz_read_value_1 = reg_file_9;
      5'b01010 : _zz_read_value_1 = reg_file_10;
      5'b01011 : _zz_read_value_1 = reg_file_11;
      5'b01100 : _zz_read_value_1 = reg_file_12;
      5'b01101 : _zz_read_value_1 = reg_file_13;
      5'b01110 : _zz_read_value_1 = reg_file_14;
      5'b01111 : _zz_read_value_1 = reg_file_15;
      5'b10000 : _zz_read_value_1 = reg_file_16;
      5'b10001 : _zz_read_value_1 = reg_file_17;
      5'b10010 : _zz_read_value_1 = reg_file_18;
      5'b10011 : _zz_read_value_1 = reg_file_19;
      5'b10100 : _zz_read_value_1 = reg_file_20;
      5'b10101 : _zz_read_value_1 = reg_file_21;
      5'b10110 : _zz_read_value_1 = reg_file_22;
      5'b10111 : _zz_read_value_1 = reg_file_23;
      5'b11000 : _zz_read_value_1 = reg_file_24;
      5'b11001 : _zz_read_value_1 = reg_file_25;
      5'b11010 : _zz_read_value_1 = reg_file_26;
      5'b11011 : _zz_read_value_1 = reg_file_27;
      5'b11100 : _zz_read_value_1 = reg_file_28;
      5'b11101 : _zz_read_value_1 = reg_file_29;
      5'b11110 : _zz_read_value_1 = reg_file_30;
      default : _zz_read_value_1 = reg_file_31;
    endcase
  end

  always @(*) begin
    case(read_ports_rs2_addr)
      5'b00000 : _zz_read_value_2 = reg_file_0;
      5'b00001 : _zz_read_value_2 = reg_file_1;
      5'b00010 : _zz_read_value_2 = reg_file_2;
      5'b00011 : _zz_read_value_2 = reg_file_3;
      5'b00100 : _zz_read_value_2 = reg_file_4;
      5'b00101 : _zz_read_value_2 = reg_file_5;
      5'b00110 : _zz_read_value_2 = reg_file_6;
      5'b00111 : _zz_read_value_2 = reg_file_7;
      5'b01000 : _zz_read_value_2 = reg_file_8;
      5'b01001 : _zz_read_value_2 = reg_file_9;
      5'b01010 : _zz_read_value_2 = reg_file_10;
      5'b01011 : _zz_read_value_2 = reg_file_11;
      5'b01100 : _zz_read_value_2 = reg_file_12;
      5'b01101 : _zz_read_value_2 = reg_file_13;
      5'b01110 : _zz_read_value_2 = reg_file_14;
      5'b01111 : _zz_read_value_2 = reg_file_15;
      5'b10000 : _zz_read_value_2 = reg_file_16;
      5'b10001 : _zz_read_value_2 = reg_file_17;
      5'b10010 : _zz_read_value_2 = reg_file_18;
      5'b10011 : _zz_read_value_2 = reg_file_19;
      5'b10100 : _zz_read_value_2 = reg_file_20;
      5'b10101 : _zz_read_value_2 = reg_file_21;
      5'b10110 : _zz_read_value_2 = reg_file_22;
      5'b10111 : _zz_read_value_2 = reg_file_23;
      5'b11000 : _zz_read_value_2 = reg_file_24;
      5'b11001 : _zz_read_value_2 = reg_file_25;
      5'b11010 : _zz_read_value_2 = reg_file_26;
      5'b11011 : _zz_read_value_2 = reg_file_27;
      5'b11100 : _zz_read_value_2 = reg_file_28;
      5'b11101 : _zz_read_value_2 = reg_file_29;
      5'b11110 : _zz_read_value_2 = reg_file_30;
      default : _zz_read_value_2 = reg_file_31;
    endcase
  end

  assign read_value_1 = _zz_read_value_1;
  assign read_value_2 = _zz_read_value_2;
  assign when_DecodePlugin_l61 = (write_ports_rd_wen && (write_ports_rd_addr != 5'h0));
  assign _zz_1 = ({31'd0,1'b1} <<< write_ports_rd_addr);
  assign read_ports_rs1_value = (((write_ports_rd_wen && ((write_ports_rd_addr == read_ports_rs1_addr) && (write_ports_rd_addr != 5'h0))) && read_ports_rs1_req) ? write_ports_rd_value : read_value_1);
  assign read_ports_rs2_value = (((write_ports_rd_wen && ((write_ports_rd_addr == read_ports_rs2_addr) && (write_ports_rd_addr != 5'h0))) && read_ports_rs2_req) ? write_ports_rd_value : read_value_2);
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      reg_file_0 <= 64'h0;
      reg_file_1 <= 64'h0;
      reg_file_2 <= 64'h0;
      reg_file_3 <= 64'h0;
      reg_file_4 <= 64'h0;
      reg_file_5 <= 64'h0;
      reg_file_6 <= 64'h0;
      reg_file_7 <= 64'h0;
      reg_file_8 <= 64'h0;
      reg_file_9 <= 64'h0;
      reg_file_10 <= 64'h0;
      reg_file_11 <= 64'h0;
      reg_file_12 <= 64'h0;
      reg_file_13 <= 64'h0;
      reg_file_14 <= 64'h0;
      reg_file_15 <= 64'h0;
      reg_file_16 <= 64'h0;
      reg_file_17 <= 64'h0;
      reg_file_18 <= 64'h0;
      reg_file_19 <= 64'h0;
      reg_file_20 <= 64'h0;
      reg_file_21 <= 64'h0;
      reg_file_22 <= 64'h0;
      reg_file_23 <= 64'h0;
      reg_file_24 <= 64'h0;
      reg_file_25 <= 64'h0;
      reg_file_26 <= 64'h0;
      reg_file_27 <= 64'h0;
      reg_file_28 <= 64'h0;
      reg_file_29 <= 64'h0;
      reg_file_30 <= 64'h0;
      reg_file_31 <= 64'h0;
    end else begin
      if(when_DecodePlugin_l61) begin
        if(_zz_1[0]) begin
          reg_file_0 <= write_ports_rd_value;
        end
        if(_zz_1[1]) begin
          reg_file_1 <= write_ports_rd_value;
        end
        if(_zz_1[2]) begin
          reg_file_2 <= write_ports_rd_value;
        end
        if(_zz_1[3]) begin
          reg_file_3 <= write_ports_rd_value;
        end
        if(_zz_1[4]) begin
          reg_file_4 <= write_ports_rd_value;
        end
        if(_zz_1[5]) begin
          reg_file_5 <= write_ports_rd_value;
        end
        if(_zz_1[6]) begin
          reg_file_6 <= write_ports_rd_value;
        end
        if(_zz_1[7]) begin
          reg_file_7 <= write_ports_rd_value;
        end
        if(_zz_1[8]) begin
          reg_file_8 <= write_ports_rd_value;
        end
        if(_zz_1[9]) begin
          reg_file_9 <= write_ports_rd_value;
        end
        if(_zz_1[10]) begin
          reg_file_10 <= write_ports_rd_value;
        end
        if(_zz_1[11]) begin
          reg_file_11 <= write_ports_rd_value;
        end
        if(_zz_1[12]) begin
          reg_file_12 <= write_ports_rd_value;
        end
        if(_zz_1[13]) begin
          reg_file_13 <= write_ports_rd_value;
        end
        if(_zz_1[14]) begin
          reg_file_14 <= write_ports_rd_value;
        end
        if(_zz_1[15]) begin
          reg_file_15 <= write_ports_rd_value;
        end
        if(_zz_1[16]) begin
          reg_file_16 <= write_ports_rd_value;
        end
        if(_zz_1[17]) begin
          reg_file_17 <= write_ports_rd_value;
        end
        if(_zz_1[18]) begin
          reg_file_18 <= write_ports_rd_value;
        end
        if(_zz_1[19]) begin
          reg_file_19 <= write_ports_rd_value;
        end
        if(_zz_1[20]) begin
          reg_file_20 <= write_ports_rd_value;
        end
        if(_zz_1[21]) begin
          reg_file_21 <= write_ports_rd_value;
        end
        if(_zz_1[22]) begin
          reg_file_22 <= write_ports_rd_value;
        end
        if(_zz_1[23]) begin
          reg_file_23 <= write_ports_rd_value;
        end
        if(_zz_1[24]) begin
          reg_file_24 <= write_ports_rd_value;
        end
        if(_zz_1[25]) begin
          reg_file_25 <= write_ports_rd_value;
        end
        if(_zz_1[26]) begin
          reg_file_26 <= write_ports_rd_value;
        end
        if(_zz_1[27]) begin
          reg_file_27 <= write_ports_rd_value;
        end
        if(_zz_1[28]) begin
          reg_file_28 <= write_ports_rd_value;
        end
        if(_zz_1[29]) begin
          reg_file_29 <= write_ports_rd_value;
        end
        if(_zz_1[30]) begin
          reg_file_30 <= write_ports_rd_value;
        end
        if(_zz_1[31]) begin
          reg_file_31 <= write_ports_rd_value;
        end
      end
    end
  end


endmodule

module gshare_predictor (
  input      [63:0]   predict_pc,
  input               predict_valid,
  output              predict_taken,
  output     [6:0]    predict_history,
  output     [63:0]   predict_pc_next,
  input               train_valid,
  input               train_taken,
  input               train_mispredicted,
  input      [6:0]    train_history,
  input      [63:0]   train_pc,
  input      [63:0]   train_pc_next,
  input               train_is_call,
  input               train_is_ret,
  input               train_is_jmp,
  input               clk,
  input               reset
);

  reg        [1:0]    _zz_GSHARE_pht_predict_taken;
  reg        [1:0]    _zz_switch_Predictor_l38;
  wire       [1:0]    _zz_BTB_btb_alloc_index_valueNext;
  wire       [0:0]    _zz_BTB_btb_alloc_index_valueNext_1;
  reg        [63:0]   _zz_RAS_ras_predict_pc;
  wire       [63:0]   _zz_predict_pc_next;
  reg        [6:0]    GSHARE_global_branch_history;
  reg        [1:0]    GSHARE_PHT_0;
  reg        [1:0]    GSHARE_PHT_1;
  reg        [1:0]    GSHARE_PHT_2;
  reg        [1:0]    GSHARE_PHT_3;
  reg        [1:0]    GSHARE_PHT_4;
  reg        [1:0]    GSHARE_PHT_5;
  reg        [1:0]    GSHARE_PHT_6;
  reg        [1:0]    GSHARE_PHT_7;
  reg        [1:0]    GSHARE_PHT_8;
  reg        [1:0]    GSHARE_PHT_9;
  reg        [1:0]    GSHARE_PHT_10;
  reg        [1:0]    GSHARE_PHT_11;
  reg        [1:0]    GSHARE_PHT_12;
  reg        [1:0]    GSHARE_PHT_13;
  reg        [1:0]    GSHARE_PHT_14;
  reg        [1:0]    GSHARE_PHT_15;
  reg        [1:0]    GSHARE_PHT_16;
  reg        [1:0]    GSHARE_PHT_17;
  reg        [1:0]    GSHARE_PHT_18;
  reg        [1:0]    GSHARE_PHT_19;
  reg        [1:0]    GSHARE_PHT_20;
  reg        [1:0]    GSHARE_PHT_21;
  reg        [1:0]    GSHARE_PHT_22;
  reg        [1:0]    GSHARE_PHT_23;
  reg        [1:0]    GSHARE_PHT_24;
  reg        [1:0]    GSHARE_PHT_25;
  reg        [1:0]    GSHARE_PHT_26;
  reg        [1:0]    GSHARE_PHT_27;
  reg        [1:0]    GSHARE_PHT_28;
  reg        [1:0]    GSHARE_PHT_29;
  reg        [1:0]    GSHARE_PHT_30;
  reg        [1:0]    GSHARE_PHT_31;
  reg        [1:0]    GSHARE_PHT_32;
  reg        [1:0]    GSHARE_PHT_33;
  reg        [1:0]    GSHARE_PHT_34;
  reg        [1:0]    GSHARE_PHT_35;
  reg        [1:0]    GSHARE_PHT_36;
  reg        [1:0]    GSHARE_PHT_37;
  reg        [1:0]    GSHARE_PHT_38;
  reg        [1:0]    GSHARE_PHT_39;
  reg        [1:0]    GSHARE_PHT_40;
  reg        [1:0]    GSHARE_PHT_41;
  reg        [1:0]    GSHARE_PHT_42;
  reg        [1:0]    GSHARE_PHT_43;
  reg        [1:0]    GSHARE_PHT_44;
  reg        [1:0]    GSHARE_PHT_45;
  reg        [1:0]    GSHARE_PHT_46;
  reg        [1:0]    GSHARE_PHT_47;
  reg        [1:0]    GSHARE_PHT_48;
  reg        [1:0]    GSHARE_PHT_49;
  reg        [1:0]    GSHARE_PHT_50;
  reg        [1:0]    GSHARE_PHT_51;
  reg        [1:0]    GSHARE_PHT_52;
  reg        [1:0]    GSHARE_PHT_53;
  reg        [1:0]    GSHARE_PHT_54;
  reg        [1:0]    GSHARE_PHT_55;
  reg        [1:0]    GSHARE_PHT_56;
  reg        [1:0]    GSHARE_PHT_57;
  reg        [1:0]    GSHARE_PHT_58;
  reg        [1:0]    GSHARE_PHT_59;
  reg        [1:0]    GSHARE_PHT_60;
  reg        [1:0]    GSHARE_PHT_61;
  reg        [1:0]    GSHARE_PHT_62;
  reg        [1:0]    GSHARE_PHT_63;
  reg        [1:0]    GSHARE_PHT_64;
  reg        [1:0]    GSHARE_PHT_65;
  reg        [1:0]    GSHARE_PHT_66;
  reg        [1:0]    GSHARE_PHT_67;
  reg        [1:0]    GSHARE_PHT_68;
  reg        [1:0]    GSHARE_PHT_69;
  reg        [1:0]    GSHARE_PHT_70;
  reg        [1:0]    GSHARE_PHT_71;
  reg        [1:0]    GSHARE_PHT_72;
  reg        [1:0]    GSHARE_PHT_73;
  reg        [1:0]    GSHARE_PHT_74;
  reg        [1:0]    GSHARE_PHT_75;
  reg        [1:0]    GSHARE_PHT_76;
  reg        [1:0]    GSHARE_PHT_77;
  reg        [1:0]    GSHARE_PHT_78;
  reg        [1:0]    GSHARE_PHT_79;
  reg        [1:0]    GSHARE_PHT_80;
  reg        [1:0]    GSHARE_PHT_81;
  reg        [1:0]    GSHARE_PHT_82;
  reg        [1:0]    GSHARE_PHT_83;
  reg        [1:0]    GSHARE_PHT_84;
  reg        [1:0]    GSHARE_PHT_85;
  reg        [1:0]    GSHARE_PHT_86;
  reg        [1:0]    GSHARE_PHT_87;
  reg        [1:0]    GSHARE_PHT_88;
  reg        [1:0]    GSHARE_PHT_89;
  reg        [1:0]    GSHARE_PHT_90;
  reg        [1:0]    GSHARE_PHT_91;
  reg        [1:0]    GSHARE_PHT_92;
  reg        [1:0]    GSHARE_PHT_93;
  reg        [1:0]    GSHARE_PHT_94;
  reg        [1:0]    GSHARE_PHT_95;
  reg        [1:0]    GSHARE_PHT_96;
  reg        [1:0]    GSHARE_PHT_97;
  reg        [1:0]    GSHARE_PHT_98;
  reg        [1:0]    GSHARE_PHT_99;
  reg        [1:0]    GSHARE_PHT_100;
  reg        [1:0]    GSHARE_PHT_101;
  reg        [1:0]    GSHARE_PHT_102;
  reg        [1:0]    GSHARE_PHT_103;
  reg        [1:0]    GSHARE_PHT_104;
  reg        [1:0]    GSHARE_PHT_105;
  reg        [1:0]    GSHARE_PHT_106;
  reg        [1:0]    GSHARE_PHT_107;
  reg        [1:0]    GSHARE_PHT_108;
  reg        [1:0]    GSHARE_PHT_109;
  reg        [1:0]    GSHARE_PHT_110;
  reg        [1:0]    GSHARE_PHT_111;
  reg        [1:0]    GSHARE_PHT_112;
  reg        [1:0]    GSHARE_PHT_113;
  reg        [1:0]    GSHARE_PHT_114;
  reg        [1:0]    GSHARE_PHT_115;
  reg        [1:0]    GSHARE_PHT_116;
  reg        [1:0]    GSHARE_PHT_117;
  reg        [1:0]    GSHARE_PHT_118;
  reg        [1:0]    GSHARE_PHT_119;
  reg        [1:0]    GSHARE_PHT_120;
  reg        [1:0]    GSHARE_PHT_121;
  reg        [1:0]    GSHARE_PHT_122;
  reg        [1:0]    GSHARE_PHT_123;
  reg        [1:0]    GSHARE_PHT_124;
  reg        [1:0]    GSHARE_PHT_125;
  reg        [1:0]    GSHARE_PHT_126;
  reg        [1:0]    GSHARE_PHT_127;
  wire       [6:0]    GSHARE_predict_index;
  wire       [6:0]    GSHARE_train_index;
  wire                GSHARE_pht_predict_taken;
  wire       [1:0]    switch_Predictor_l38;
  wire       [127:0]  _zz_1;
  wire                _zz_2;
  wire                _zz_3;
  wire                _zz_4;
  wire                _zz_5;
  wire                _zz_6;
  wire                _zz_7;
  wire                _zz_8;
  wire                _zz_9;
  wire                _zz_10;
  wire                _zz_11;
  wire                _zz_12;
  wire                _zz_13;
  wire                _zz_14;
  wire                _zz_15;
  wire                _zz_16;
  wire                _zz_17;
  wire                _zz_18;
  wire                _zz_19;
  wire                _zz_20;
  wire                _zz_21;
  wire                _zz_22;
  wire                _zz_23;
  wire                _zz_24;
  wire                _zz_25;
  wire                _zz_26;
  wire                _zz_27;
  wire                _zz_28;
  wire                _zz_29;
  wire                _zz_30;
  wire                _zz_31;
  wire                _zz_32;
  wire                _zz_33;
  wire                _zz_34;
  wire                _zz_35;
  wire                _zz_36;
  wire                _zz_37;
  wire                _zz_38;
  wire                _zz_39;
  wire                _zz_40;
  wire                _zz_41;
  wire                _zz_42;
  wire                _zz_43;
  wire                _zz_44;
  wire                _zz_45;
  wire                _zz_46;
  wire                _zz_47;
  wire                _zz_48;
  wire                _zz_49;
  wire                _zz_50;
  wire                _zz_51;
  wire                _zz_52;
  wire                _zz_53;
  wire                _zz_54;
  wire                _zz_55;
  wire                _zz_56;
  wire                _zz_57;
  wire                _zz_58;
  wire                _zz_59;
  wire                _zz_60;
  wire                _zz_61;
  wire                _zz_62;
  wire                _zz_63;
  wire                _zz_64;
  wire                _zz_65;
  wire                _zz_66;
  wire                _zz_67;
  wire                _zz_68;
  wire                _zz_69;
  wire                _zz_70;
  wire                _zz_71;
  wire                _zz_72;
  wire                _zz_73;
  wire                _zz_74;
  wire                _zz_75;
  wire                _zz_76;
  wire                _zz_77;
  wire                _zz_78;
  wire                _zz_79;
  wire                _zz_80;
  wire                _zz_81;
  wire                _zz_82;
  wire                _zz_83;
  wire                _zz_84;
  wire                _zz_85;
  wire                _zz_86;
  wire                _zz_87;
  wire                _zz_88;
  wire                _zz_89;
  wire                _zz_90;
  wire                _zz_91;
  wire                _zz_92;
  wire                _zz_93;
  wire                _zz_94;
  wire                _zz_95;
  wire                _zz_96;
  wire                _zz_97;
  wire                _zz_98;
  wire                _zz_99;
  wire                _zz_100;
  wire                _zz_101;
  wire                _zz_102;
  wire                _zz_103;
  wire                _zz_104;
  wire                _zz_105;
  wire                _zz_106;
  wire                _zz_107;
  wire                _zz_108;
  wire                _zz_109;
  wire                _zz_110;
  wire                _zz_111;
  wire                _zz_112;
  wire                _zz_113;
  wire                _zz_114;
  wire                _zz_115;
  wire                _zz_116;
  wire                _zz_117;
  wire                _zz_118;
  wire                _zz_119;
  wire                _zz_120;
  wire                _zz_121;
  wire                _zz_122;
  wire                _zz_123;
  wire                _zz_124;
  wire                _zz_125;
  wire                _zz_126;
  wire                _zz_127;
  wire                _zz_128;
  wire                _zz_129;
  wire                when_Predictor_l61;
  wire                when_Predictor_l70;
  reg        [3:0]    BTB_valid;
  reg        [63:0]   BTB_source_pc_0;
  reg        [63:0]   BTB_source_pc_1;
  reg        [63:0]   BTB_source_pc_2;
  reg        [63:0]   BTB_source_pc_3;
  reg        [3:0]    BTB_call;
  reg        [3:0]    BTB_ret;
  reg        [3:0]    BTB_jmp;
  reg        [63:0]   BTB_target_pc_0;
  reg        [63:0]   BTB_target_pc_1;
  reg        [63:0]   BTB_target_pc_2;
  reg        [63:0]   BTB_target_pc_3;
  reg                 BTB_is_matched;
  reg                 BTB_is_call;
  reg                 BTB_is_ret;
  reg                 BTB_is_jmp;
  reg        [63:0]   BTB_target_pc_read;
  wire                when_Predictor_l95;
  wire                when_Predictor_l95_1;
  wire                when_Predictor_l95_2;
  wire                when_Predictor_l95_3;
  wire       [1:0]    BTB_btb_write_index;
  reg                 BTB_btb_alloc_index_willIncrement;
  reg                 BTB_btb_alloc_index_willClear;
  reg        [1:0]    BTB_btb_alloc_index_valueNext;
  reg        [1:0]    BTB_btb_alloc_index_value;
  wire                BTB_btb_alloc_index_willOverflowIfInc;
  wire                BTB_btb_alloc_index_willOverflow;
  reg                 BTB_btb_is_hit_vec_0;
  reg                 BTB_btb_is_hit_vec_1;
  reg                 BTB_btb_is_hit_vec_2;
  reg                 BTB_btb_is_hit_vec_3;
  reg                 BTB_btb_is_miss_vec_0;
  reg                 BTB_btb_is_miss_vec_1;
  reg                 BTB_btb_is_miss_vec_2;
  reg                 BTB_btb_is_miss_vec_3;
  wire                BTB_btb_is_hit;
  wire                BTB_btb_is_miss;
  wire                when_Predictor_l113;
  wire                when_Predictor_l114;
  wire                when_Predictor_l119;
  wire                when_Predictor_l113_1;
  wire                when_Predictor_l114_1;
  wire                when_Predictor_l119_1;
  wire                when_Predictor_l113_2;
  wire                when_Predictor_l114_2;
  wire                when_Predictor_l119_2;
  wire                when_Predictor_l113_3;
  wire                when_Predictor_l114_3;
  wire                when_Predictor_l119_3;
  wire                _zz_BTB_btb_write_index;
  wire                _zz_BTB_btb_write_index_1;
  wire       [3:0]    _zz_130;
  wire       [3:0]    _zz_131;
  wire       [3:0]    _zz_132;
  wire       [3:0]    _zz_133;
  reg        [63:0]   RAS_ras_regfile_0;
  reg        [63:0]   RAS_ras_regfile_1;
  reg        [63:0]   RAS_ras_regfile_2;
  reg        [63:0]   RAS_ras_regfile_3;
  reg        [1:0]    RAS_ras_next_index;
  reg        [1:0]    RAS_ras_curr_index;
  reg        [1:0]    RAS_ras_next_index_proven;
  reg        [1:0]    RAS_ras_curr_index_proven;
  wire       [63:0]   RAS_ras_predict_pc;
  wire                RAS_ras_call_matched;
  wire                RAS_ras_ret_matched;
  wire                when_Predictor_l169;
  wire                when_Predictor_l172;
  wire                when_Predictor_l180;
  wire                when_Predictor_l183;
  wire                when_Predictor_l197;
  wire       [3:0]    _zz_134;
  wire                _zz_135;
  wire                _zz_136;
  wire                _zz_137;
  wire                _zz_138;
  wire       [63:0]   _zz_RAS_ras_regfile_0;
  wire       [63:0]   _zz_RAS_ras_regfile_0_1;
  wire                when_Predictor_l205;

  assign _zz_BTB_btb_alloc_index_valueNext_1 = BTB_btb_alloc_index_willIncrement;
  assign _zz_BTB_btb_alloc_index_valueNext = {1'd0, _zz_BTB_btb_alloc_index_valueNext_1};
  assign _zz_predict_pc_next = (predict_pc + 64'h0000000000000004);
  always @(*) begin
    case(GSHARE_predict_index)
      7'b0000000 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_0;
      7'b0000001 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_1;
      7'b0000010 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_2;
      7'b0000011 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_3;
      7'b0000100 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_4;
      7'b0000101 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_5;
      7'b0000110 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_6;
      7'b0000111 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_7;
      7'b0001000 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_8;
      7'b0001001 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_9;
      7'b0001010 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_10;
      7'b0001011 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_11;
      7'b0001100 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_12;
      7'b0001101 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_13;
      7'b0001110 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_14;
      7'b0001111 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_15;
      7'b0010000 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_16;
      7'b0010001 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_17;
      7'b0010010 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_18;
      7'b0010011 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_19;
      7'b0010100 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_20;
      7'b0010101 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_21;
      7'b0010110 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_22;
      7'b0010111 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_23;
      7'b0011000 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_24;
      7'b0011001 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_25;
      7'b0011010 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_26;
      7'b0011011 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_27;
      7'b0011100 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_28;
      7'b0011101 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_29;
      7'b0011110 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_30;
      7'b0011111 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_31;
      7'b0100000 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_32;
      7'b0100001 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_33;
      7'b0100010 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_34;
      7'b0100011 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_35;
      7'b0100100 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_36;
      7'b0100101 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_37;
      7'b0100110 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_38;
      7'b0100111 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_39;
      7'b0101000 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_40;
      7'b0101001 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_41;
      7'b0101010 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_42;
      7'b0101011 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_43;
      7'b0101100 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_44;
      7'b0101101 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_45;
      7'b0101110 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_46;
      7'b0101111 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_47;
      7'b0110000 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_48;
      7'b0110001 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_49;
      7'b0110010 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_50;
      7'b0110011 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_51;
      7'b0110100 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_52;
      7'b0110101 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_53;
      7'b0110110 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_54;
      7'b0110111 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_55;
      7'b0111000 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_56;
      7'b0111001 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_57;
      7'b0111010 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_58;
      7'b0111011 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_59;
      7'b0111100 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_60;
      7'b0111101 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_61;
      7'b0111110 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_62;
      7'b0111111 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_63;
      7'b1000000 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_64;
      7'b1000001 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_65;
      7'b1000010 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_66;
      7'b1000011 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_67;
      7'b1000100 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_68;
      7'b1000101 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_69;
      7'b1000110 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_70;
      7'b1000111 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_71;
      7'b1001000 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_72;
      7'b1001001 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_73;
      7'b1001010 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_74;
      7'b1001011 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_75;
      7'b1001100 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_76;
      7'b1001101 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_77;
      7'b1001110 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_78;
      7'b1001111 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_79;
      7'b1010000 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_80;
      7'b1010001 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_81;
      7'b1010010 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_82;
      7'b1010011 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_83;
      7'b1010100 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_84;
      7'b1010101 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_85;
      7'b1010110 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_86;
      7'b1010111 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_87;
      7'b1011000 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_88;
      7'b1011001 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_89;
      7'b1011010 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_90;
      7'b1011011 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_91;
      7'b1011100 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_92;
      7'b1011101 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_93;
      7'b1011110 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_94;
      7'b1011111 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_95;
      7'b1100000 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_96;
      7'b1100001 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_97;
      7'b1100010 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_98;
      7'b1100011 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_99;
      7'b1100100 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_100;
      7'b1100101 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_101;
      7'b1100110 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_102;
      7'b1100111 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_103;
      7'b1101000 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_104;
      7'b1101001 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_105;
      7'b1101010 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_106;
      7'b1101011 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_107;
      7'b1101100 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_108;
      7'b1101101 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_109;
      7'b1101110 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_110;
      7'b1101111 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_111;
      7'b1110000 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_112;
      7'b1110001 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_113;
      7'b1110010 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_114;
      7'b1110011 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_115;
      7'b1110100 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_116;
      7'b1110101 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_117;
      7'b1110110 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_118;
      7'b1110111 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_119;
      7'b1111000 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_120;
      7'b1111001 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_121;
      7'b1111010 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_122;
      7'b1111011 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_123;
      7'b1111100 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_124;
      7'b1111101 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_125;
      7'b1111110 : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_126;
      default : _zz_GSHARE_pht_predict_taken = GSHARE_PHT_127;
    endcase
  end

  always @(*) begin
    case(GSHARE_train_index)
      7'b0000000 : _zz_switch_Predictor_l38 = GSHARE_PHT_0;
      7'b0000001 : _zz_switch_Predictor_l38 = GSHARE_PHT_1;
      7'b0000010 : _zz_switch_Predictor_l38 = GSHARE_PHT_2;
      7'b0000011 : _zz_switch_Predictor_l38 = GSHARE_PHT_3;
      7'b0000100 : _zz_switch_Predictor_l38 = GSHARE_PHT_4;
      7'b0000101 : _zz_switch_Predictor_l38 = GSHARE_PHT_5;
      7'b0000110 : _zz_switch_Predictor_l38 = GSHARE_PHT_6;
      7'b0000111 : _zz_switch_Predictor_l38 = GSHARE_PHT_7;
      7'b0001000 : _zz_switch_Predictor_l38 = GSHARE_PHT_8;
      7'b0001001 : _zz_switch_Predictor_l38 = GSHARE_PHT_9;
      7'b0001010 : _zz_switch_Predictor_l38 = GSHARE_PHT_10;
      7'b0001011 : _zz_switch_Predictor_l38 = GSHARE_PHT_11;
      7'b0001100 : _zz_switch_Predictor_l38 = GSHARE_PHT_12;
      7'b0001101 : _zz_switch_Predictor_l38 = GSHARE_PHT_13;
      7'b0001110 : _zz_switch_Predictor_l38 = GSHARE_PHT_14;
      7'b0001111 : _zz_switch_Predictor_l38 = GSHARE_PHT_15;
      7'b0010000 : _zz_switch_Predictor_l38 = GSHARE_PHT_16;
      7'b0010001 : _zz_switch_Predictor_l38 = GSHARE_PHT_17;
      7'b0010010 : _zz_switch_Predictor_l38 = GSHARE_PHT_18;
      7'b0010011 : _zz_switch_Predictor_l38 = GSHARE_PHT_19;
      7'b0010100 : _zz_switch_Predictor_l38 = GSHARE_PHT_20;
      7'b0010101 : _zz_switch_Predictor_l38 = GSHARE_PHT_21;
      7'b0010110 : _zz_switch_Predictor_l38 = GSHARE_PHT_22;
      7'b0010111 : _zz_switch_Predictor_l38 = GSHARE_PHT_23;
      7'b0011000 : _zz_switch_Predictor_l38 = GSHARE_PHT_24;
      7'b0011001 : _zz_switch_Predictor_l38 = GSHARE_PHT_25;
      7'b0011010 : _zz_switch_Predictor_l38 = GSHARE_PHT_26;
      7'b0011011 : _zz_switch_Predictor_l38 = GSHARE_PHT_27;
      7'b0011100 : _zz_switch_Predictor_l38 = GSHARE_PHT_28;
      7'b0011101 : _zz_switch_Predictor_l38 = GSHARE_PHT_29;
      7'b0011110 : _zz_switch_Predictor_l38 = GSHARE_PHT_30;
      7'b0011111 : _zz_switch_Predictor_l38 = GSHARE_PHT_31;
      7'b0100000 : _zz_switch_Predictor_l38 = GSHARE_PHT_32;
      7'b0100001 : _zz_switch_Predictor_l38 = GSHARE_PHT_33;
      7'b0100010 : _zz_switch_Predictor_l38 = GSHARE_PHT_34;
      7'b0100011 : _zz_switch_Predictor_l38 = GSHARE_PHT_35;
      7'b0100100 : _zz_switch_Predictor_l38 = GSHARE_PHT_36;
      7'b0100101 : _zz_switch_Predictor_l38 = GSHARE_PHT_37;
      7'b0100110 : _zz_switch_Predictor_l38 = GSHARE_PHT_38;
      7'b0100111 : _zz_switch_Predictor_l38 = GSHARE_PHT_39;
      7'b0101000 : _zz_switch_Predictor_l38 = GSHARE_PHT_40;
      7'b0101001 : _zz_switch_Predictor_l38 = GSHARE_PHT_41;
      7'b0101010 : _zz_switch_Predictor_l38 = GSHARE_PHT_42;
      7'b0101011 : _zz_switch_Predictor_l38 = GSHARE_PHT_43;
      7'b0101100 : _zz_switch_Predictor_l38 = GSHARE_PHT_44;
      7'b0101101 : _zz_switch_Predictor_l38 = GSHARE_PHT_45;
      7'b0101110 : _zz_switch_Predictor_l38 = GSHARE_PHT_46;
      7'b0101111 : _zz_switch_Predictor_l38 = GSHARE_PHT_47;
      7'b0110000 : _zz_switch_Predictor_l38 = GSHARE_PHT_48;
      7'b0110001 : _zz_switch_Predictor_l38 = GSHARE_PHT_49;
      7'b0110010 : _zz_switch_Predictor_l38 = GSHARE_PHT_50;
      7'b0110011 : _zz_switch_Predictor_l38 = GSHARE_PHT_51;
      7'b0110100 : _zz_switch_Predictor_l38 = GSHARE_PHT_52;
      7'b0110101 : _zz_switch_Predictor_l38 = GSHARE_PHT_53;
      7'b0110110 : _zz_switch_Predictor_l38 = GSHARE_PHT_54;
      7'b0110111 : _zz_switch_Predictor_l38 = GSHARE_PHT_55;
      7'b0111000 : _zz_switch_Predictor_l38 = GSHARE_PHT_56;
      7'b0111001 : _zz_switch_Predictor_l38 = GSHARE_PHT_57;
      7'b0111010 : _zz_switch_Predictor_l38 = GSHARE_PHT_58;
      7'b0111011 : _zz_switch_Predictor_l38 = GSHARE_PHT_59;
      7'b0111100 : _zz_switch_Predictor_l38 = GSHARE_PHT_60;
      7'b0111101 : _zz_switch_Predictor_l38 = GSHARE_PHT_61;
      7'b0111110 : _zz_switch_Predictor_l38 = GSHARE_PHT_62;
      7'b0111111 : _zz_switch_Predictor_l38 = GSHARE_PHT_63;
      7'b1000000 : _zz_switch_Predictor_l38 = GSHARE_PHT_64;
      7'b1000001 : _zz_switch_Predictor_l38 = GSHARE_PHT_65;
      7'b1000010 : _zz_switch_Predictor_l38 = GSHARE_PHT_66;
      7'b1000011 : _zz_switch_Predictor_l38 = GSHARE_PHT_67;
      7'b1000100 : _zz_switch_Predictor_l38 = GSHARE_PHT_68;
      7'b1000101 : _zz_switch_Predictor_l38 = GSHARE_PHT_69;
      7'b1000110 : _zz_switch_Predictor_l38 = GSHARE_PHT_70;
      7'b1000111 : _zz_switch_Predictor_l38 = GSHARE_PHT_71;
      7'b1001000 : _zz_switch_Predictor_l38 = GSHARE_PHT_72;
      7'b1001001 : _zz_switch_Predictor_l38 = GSHARE_PHT_73;
      7'b1001010 : _zz_switch_Predictor_l38 = GSHARE_PHT_74;
      7'b1001011 : _zz_switch_Predictor_l38 = GSHARE_PHT_75;
      7'b1001100 : _zz_switch_Predictor_l38 = GSHARE_PHT_76;
      7'b1001101 : _zz_switch_Predictor_l38 = GSHARE_PHT_77;
      7'b1001110 : _zz_switch_Predictor_l38 = GSHARE_PHT_78;
      7'b1001111 : _zz_switch_Predictor_l38 = GSHARE_PHT_79;
      7'b1010000 : _zz_switch_Predictor_l38 = GSHARE_PHT_80;
      7'b1010001 : _zz_switch_Predictor_l38 = GSHARE_PHT_81;
      7'b1010010 : _zz_switch_Predictor_l38 = GSHARE_PHT_82;
      7'b1010011 : _zz_switch_Predictor_l38 = GSHARE_PHT_83;
      7'b1010100 : _zz_switch_Predictor_l38 = GSHARE_PHT_84;
      7'b1010101 : _zz_switch_Predictor_l38 = GSHARE_PHT_85;
      7'b1010110 : _zz_switch_Predictor_l38 = GSHARE_PHT_86;
      7'b1010111 : _zz_switch_Predictor_l38 = GSHARE_PHT_87;
      7'b1011000 : _zz_switch_Predictor_l38 = GSHARE_PHT_88;
      7'b1011001 : _zz_switch_Predictor_l38 = GSHARE_PHT_89;
      7'b1011010 : _zz_switch_Predictor_l38 = GSHARE_PHT_90;
      7'b1011011 : _zz_switch_Predictor_l38 = GSHARE_PHT_91;
      7'b1011100 : _zz_switch_Predictor_l38 = GSHARE_PHT_92;
      7'b1011101 : _zz_switch_Predictor_l38 = GSHARE_PHT_93;
      7'b1011110 : _zz_switch_Predictor_l38 = GSHARE_PHT_94;
      7'b1011111 : _zz_switch_Predictor_l38 = GSHARE_PHT_95;
      7'b1100000 : _zz_switch_Predictor_l38 = GSHARE_PHT_96;
      7'b1100001 : _zz_switch_Predictor_l38 = GSHARE_PHT_97;
      7'b1100010 : _zz_switch_Predictor_l38 = GSHARE_PHT_98;
      7'b1100011 : _zz_switch_Predictor_l38 = GSHARE_PHT_99;
      7'b1100100 : _zz_switch_Predictor_l38 = GSHARE_PHT_100;
      7'b1100101 : _zz_switch_Predictor_l38 = GSHARE_PHT_101;
      7'b1100110 : _zz_switch_Predictor_l38 = GSHARE_PHT_102;
      7'b1100111 : _zz_switch_Predictor_l38 = GSHARE_PHT_103;
      7'b1101000 : _zz_switch_Predictor_l38 = GSHARE_PHT_104;
      7'b1101001 : _zz_switch_Predictor_l38 = GSHARE_PHT_105;
      7'b1101010 : _zz_switch_Predictor_l38 = GSHARE_PHT_106;
      7'b1101011 : _zz_switch_Predictor_l38 = GSHARE_PHT_107;
      7'b1101100 : _zz_switch_Predictor_l38 = GSHARE_PHT_108;
      7'b1101101 : _zz_switch_Predictor_l38 = GSHARE_PHT_109;
      7'b1101110 : _zz_switch_Predictor_l38 = GSHARE_PHT_110;
      7'b1101111 : _zz_switch_Predictor_l38 = GSHARE_PHT_111;
      7'b1110000 : _zz_switch_Predictor_l38 = GSHARE_PHT_112;
      7'b1110001 : _zz_switch_Predictor_l38 = GSHARE_PHT_113;
      7'b1110010 : _zz_switch_Predictor_l38 = GSHARE_PHT_114;
      7'b1110011 : _zz_switch_Predictor_l38 = GSHARE_PHT_115;
      7'b1110100 : _zz_switch_Predictor_l38 = GSHARE_PHT_116;
      7'b1110101 : _zz_switch_Predictor_l38 = GSHARE_PHT_117;
      7'b1110110 : _zz_switch_Predictor_l38 = GSHARE_PHT_118;
      7'b1110111 : _zz_switch_Predictor_l38 = GSHARE_PHT_119;
      7'b1111000 : _zz_switch_Predictor_l38 = GSHARE_PHT_120;
      7'b1111001 : _zz_switch_Predictor_l38 = GSHARE_PHT_121;
      7'b1111010 : _zz_switch_Predictor_l38 = GSHARE_PHT_122;
      7'b1111011 : _zz_switch_Predictor_l38 = GSHARE_PHT_123;
      7'b1111100 : _zz_switch_Predictor_l38 = GSHARE_PHT_124;
      7'b1111101 : _zz_switch_Predictor_l38 = GSHARE_PHT_125;
      7'b1111110 : _zz_switch_Predictor_l38 = GSHARE_PHT_126;
      default : _zz_switch_Predictor_l38 = GSHARE_PHT_127;
    endcase
  end

  always @(*) begin
    case(RAS_ras_curr_index)
      2'b00 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_0;
      2'b01 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_1;
      2'b10 : _zz_RAS_ras_predict_pc = RAS_ras_regfile_2;
      default : _zz_RAS_ras_predict_pc = RAS_ras_regfile_3;
    endcase
  end

  assign GSHARE_predict_index = (predict_pc[8 : 2] ^ GSHARE_global_branch_history);
  assign GSHARE_train_index = (train_pc[8 : 2] ^ train_history);
  assign GSHARE_pht_predict_taken = _zz_GSHARE_pht_predict_taken[1];
  assign switch_Predictor_l38 = _zz_switch_Predictor_l38;
  assign _zz_1 = ({127'd0,1'b1} <<< GSHARE_train_index);
  assign _zz_2 = _zz_1[0];
  assign _zz_3 = _zz_1[1];
  assign _zz_4 = _zz_1[2];
  assign _zz_5 = _zz_1[3];
  assign _zz_6 = _zz_1[4];
  assign _zz_7 = _zz_1[5];
  assign _zz_8 = _zz_1[6];
  assign _zz_9 = _zz_1[7];
  assign _zz_10 = _zz_1[8];
  assign _zz_11 = _zz_1[9];
  assign _zz_12 = _zz_1[10];
  assign _zz_13 = _zz_1[11];
  assign _zz_14 = _zz_1[12];
  assign _zz_15 = _zz_1[13];
  assign _zz_16 = _zz_1[14];
  assign _zz_17 = _zz_1[15];
  assign _zz_18 = _zz_1[16];
  assign _zz_19 = _zz_1[17];
  assign _zz_20 = _zz_1[18];
  assign _zz_21 = _zz_1[19];
  assign _zz_22 = _zz_1[20];
  assign _zz_23 = _zz_1[21];
  assign _zz_24 = _zz_1[22];
  assign _zz_25 = _zz_1[23];
  assign _zz_26 = _zz_1[24];
  assign _zz_27 = _zz_1[25];
  assign _zz_28 = _zz_1[26];
  assign _zz_29 = _zz_1[27];
  assign _zz_30 = _zz_1[28];
  assign _zz_31 = _zz_1[29];
  assign _zz_32 = _zz_1[30];
  assign _zz_33 = _zz_1[31];
  assign _zz_34 = _zz_1[32];
  assign _zz_35 = _zz_1[33];
  assign _zz_36 = _zz_1[34];
  assign _zz_37 = _zz_1[35];
  assign _zz_38 = _zz_1[36];
  assign _zz_39 = _zz_1[37];
  assign _zz_40 = _zz_1[38];
  assign _zz_41 = _zz_1[39];
  assign _zz_42 = _zz_1[40];
  assign _zz_43 = _zz_1[41];
  assign _zz_44 = _zz_1[42];
  assign _zz_45 = _zz_1[43];
  assign _zz_46 = _zz_1[44];
  assign _zz_47 = _zz_1[45];
  assign _zz_48 = _zz_1[46];
  assign _zz_49 = _zz_1[47];
  assign _zz_50 = _zz_1[48];
  assign _zz_51 = _zz_1[49];
  assign _zz_52 = _zz_1[50];
  assign _zz_53 = _zz_1[51];
  assign _zz_54 = _zz_1[52];
  assign _zz_55 = _zz_1[53];
  assign _zz_56 = _zz_1[54];
  assign _zz_57 = _zz_1[55];
  assign _zz_58 = _zz_1[56];
  assign _zz_59 = _zz_1[57];
  assign _zz_60 = _zz_1[58];
  assign _zz_61 = _zz_1[59];
  assign _zz_62 = _zz_1[60];
  assign _zz_63 = _zz_1[61];
  assign _zz_64 = _zz_1[62];
  assign _zz_65 = _zz_1[63];
  assign _zz_66 = _zz_1[64];
  assign _zz_67 = _zz_1[65];
  assign _zz_68 = _zz_1[66];
  assign _zz_69 = _zz_1[67];
  assign _zz_70 = _zz_1[68];
  assign _zz_71 = _zz_1[69];
  assign _zz_72 = _zz_1[70];
  assign _zz_73 = _zz_1[71];
  assign _zz_74 = _zz_1[72];
  assign _zz_75 = _zz_1[73];
  assign _zz_76 = _zz_1[74];
  assign _zz_77 = _zz_1[75];
  assign _zz_78 = _zz_1[76];
  assign _zz_79 = _zz_1[77];
  assign _zz_80 = _zz_1[78];
  assign _zz_81 = _zz_1[79];
  assign _zz_82 = _zz_1[80];
  assign _zz_83 = _zz_1[81];
  assign _zz_84 = _zz_1[82];
  assign _zz_85 = _zz_1[83];
  assign _zz_86 = _zz_1[84];
  assign _zz_87 = _zz_1[85];
  assign _zz_88 = _zz_1[86];
  assign _zz_89 = _zz_1[87];
  assign _zz_90 = _zz_1[88];
  assign _zz_91 = _zz_1[89];
  assign _zz_92 = _zz_1[90];
  assign _zz_93 = _zz_1[91];
  assign _zz_94 = _zz_1[92];
  assign _zz_95 = _zz_1[93];
  assign _zz_96 = _zz_1[94];
  assign _zz_97 = _zz_1[95];
  assign _zz_98 = _zz_1[96];
  assign _zz_99 = _zz_1[97];
  assign _zz_100 = _zz_1[98];
  assign _zz_101 = _zz_1[99];
  assign _zz_102 = _zz_1[100];
  assign _zz_103 = _zz_1[101];
  assign _zz_104 = _zz_1[102];
  assign _zz_105 = _zz_1[103];
  assign _zz_106 = _zz_1[104];
  assign _zz_107 = _zz_1[105];
  assign _zz_108 = _zz_1[106];
  assign _zz_109 = _zz_1[107];
  assign _zz_110 = _zz_1[108];
  assign _zz_111 = _zz_1[109];
  assign _zz_112 = _zz_1[110];
  assign _zz_113 = _zz_1[111];
  assign _zz_114 = _zz_1[112];
  assign _zz_115 = _zz_1[113];
  assign _zz_116 = _zz_1[114];
  assign _zz_117 = _zz_1[115];
  assign _zz_118 = _zz_1[116];
  assign _zz_119 = _zz_1[117];
  assign _zz_120 = _zz_1[118];
  assign _zz_121 = _zz_1[119];
  assign _zz_122 = _zz_1[120];
  assign _zz_123 = _zz_1[121];
  assign _zz_124 = _zz_1[122];
  assign _zz_125 = _zz_1[123];
  assign _zz_126 = _zz_1[124];
  assign _zz_127 = _zz_1[125];
  assign _zz_128 = _zz_1[126];
  assign _zz_129 = _zz_1[127];
  assign when_Predictor_l61 = (! train_taken);
  assign when_Predictor_l70 = (train_valid && train_mispredicted);
  always @(*) begin
    BTB_is_matched = 1'b0;
    if(when_Predictor_l95) begin
      BTB_is_matched = 1'b1;
    end
    if(when_Predictor_l95_1) begin
      BTB_is_matched = 1'b1;
    end
    if(when_Predictor_l95_2) begin
      BTB_is_matched = 1'b1;
    end
    if(when_Predictor_l95_3) begin
      BTB_is_matched = 1'b1;
    end
  end

  always @(*) begin
    BTB_is_call = 1'b0;
    if(when_Predictor_l95) begin
      BTB_is_call = BTB_call[0];
    end
    if(when_Predictor_l95_1) begin
      BTB_is_call = BTB_call[1];
    end
    if(when_Predictor_l95_2) begin
      BTB_is_call = BTB_call[2];
    end
    if(when_Predictor_l95_3) begin
      BTB_is_call = BTB_call[3];
    end
  end

  always @(*) begin
    BTB_is_ret = 1'b0;
    if(when_Predictor_l95) begin
      BTB_is_ret = BTB_ret[0];
    end
    if(when_Predictor_l95_1) begin
      BTB_is_ret = BTB_ret[1];
    end
    if(when_Predictor_l95_2) begin
      BTB_is_ret = BTB_ret[2];
    end
    if(when_Predictor_l95_3) begin
      BTB_is_ret = BTB_ret[3];
    end
  end

  always @(*) begin
    BTB_is_jmp = 1'b0;
    if(when_Predictor_l95) begin
      BTB_is_jmp = BTB_jmp[0];
    end
    if(when_Predictor_l95_1) begin
      BTB_is_jmp = BTB_jmp[1];
    end
    if(when_Predictor_l95_2) begin
      BTB_is_jmp = BTB_jmp[2];
    end
    if(when_Predictor_l95_3) begin
      BTB_is_jmp = BTB_jmp[3];
    end
  end

  always @(*) begin
    BTB_target_pc_read = 64'h0;
    if(when_Predictor_l95) begin
      BTB_target_pc_read = BTB_target_pc_0;
    end
    if(when_Predictor_l95_1) begin
      BTB_target_pc_read = BTB_target_pc_1;
    end
    if(when_Predictor_l95_2) begin
      BTB_target_pc_read = BTB_target_pc_2;
    end
    if(when_Predictor_l95_3) begin
      BTB_target_pc_read = BTB_target_pc_3;
    end
  end

  assign when_Predictor_l95 = ((BTB_source_pc_0 == predict_pc) && BTB_valid[0]);
  assign when_Predictor_l95_1 = ((BTB_source_pc_1 == predict_pc) && BTB_valid[1]);
  assign when_Predictor_l95_2 = ((BTB_source_pc_2 == predict_pc) && BTB_valid[2]);
  assign when_Predictor_l95_3 = ((BTB_source_pc_3 == predict_pc) && BTB_valid[3]);
  always @(*) begin
    BTB_btb_alloc_index_willIncrement = 1'b0;
    if(BTB_btb_is_miss) begin
      if(!BTB_btb_alloc_index_willOverflowIfInc) begin
        BTB_btb_alloc_index_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    BTB_btb_alloc_index_willClear = 1'b0;
    if(BTB_btb_is_miss) begin
      if(BTB_btb_alloc_index_willOverflowIfInc) begin
        BTB_btb_alloc_index_willClear = 1'b1;
      end
    end
  end

  assign BTB_btb_alloc_index_willOverflowIfInc = (BTB_btb_alloc_index_value == 2'b11);
  assign BTB_btb_alloc_index_willOverflow = (BTB_btb_alloc_index_willOverflowIfInc && BTB_btb_alloc_index_willIncrement);
  always @(*) begin
    BTB_btb_alloc_index_valueNext = (BTB_btb_alloc_index_value + _zz_BTB_btb_alloc_index_valueNext);
    if(BTB_btb_alloc_index_willClear) begin
      BTB_btb_alloc_index_valueNext = 2'b00;
    end
  end

  assign BTB_btb_is_hit = (|{BTB_btb_is_hit_vec_3,{BTB_btb_is_hit_vec_2,{BTB_btb_is_hit_vec_1,BTB_btb_is_hit_vec_0}}});
  assign BTB_btb_is_miss = (|{BTB_btb_is_miss_vec_3,{BTB_btb_is_miss_vec_2,{BTB_btb_is_miss_vec_1,BTB_btb_is_miss_vec_0}}});
  assign when_Predictor_l113 = (train_valid && train_taken);
  assign when_Predictor_l114 = ((BTB_source_pc_0 == train_pc) && BTB_valid[0]);
  always @(*) begin
    if(when_Predictor_l113) begin
      if(when_Predictor_l114) begin
        BTB_btb_is_hit_vec_0 = 1'b1;
      end else begin
        BTB_btb_is_hit_vec_0 = 1'b0;
      end
    end else begin
      BTB_btb_is_hit_vec_0 = 1'b0;
    end
  end

  assign when_Predictor_l119 = ((BTB_source_pc_0 != train_pc) || (! BTB_valid[0]));
  always @(*) begin
    if(when_Predictor_l113) begin
      if(when_Predictor_l119) begin
        BTB_btb_is_miss_vec_0 = 1'b1;
      end else begin
        BTB_btb_is_miss_vec_0 = 1'b0;
      end
    end else begin
      BTB_btb_is_miss_vec_0 = 1'b0;
    end
  end

  assign when_Predictor_l113_1 = (train_valid && train_taken);
  assign when_Predictor_l114_1 = ((BTB_source_pc_1 == train_pc) && BTB_valid[1]);
  always @(*) begin
    if(when_Predictor_l113_1) begin
      if(when_Predictor_l114_1) begin
        BTB_btb_is_hit_vec_1 = 1'b1;
      end else begin
        BTB_btb_is_hit_vec_1 = 1'b0;
      end
    end else begin
      BTB_btb_is_hit_vec_1 = 1'b0;
    end
  end

  assign when_Predictor_l119_1 = ((BTB_source_pc_1 != train_pc) || (! BTB_valid[1]));
  always @(*) begin
    if(when_Predictor_l113_1) begin
      if(when_Predictor_l119_1) begin
        BTB_btb_is_miss_vec_1 = 1'b1;
      end else begin
        BTB_btb_is_miss_vec_1 = 1'b0;
      end
    end else begin
      BTB_btb_is_miss_vec_1 = 1'b0;
    end
  end

  assign when_Predictor_l113_2 = (train_valid && train_taken);
  assign when_Predictor_l114_2 = ((BTB_source_pc_2 == train_pc) && BTB_valid[2]);
  always @(*) begin
    if(when_Predictor_l113_2) begin
      if(when_Predictor_l114_2) begin
        BTB_btb_is_hit_vec_2 = 1'b1;
      end else begin
        BTB_btb_is_hit_vec_2 = 1'b0;
      end
    end else begin
      BTB_btb_is_hit_vec_2 = 1'b0;
    end
  end

  assign when_Predictor_l119_2 = ((BTB_source_pc_2 != train_pc) || (! BTB_valid[2]));
  always @(*) begin
    if(when_Predictor_l113_2) begin
      if(when_Predictor_l119_2) begin
        BTB_btb_is_miss_vec_2 = 1'b1;
      end else begin
        BTB_btb_is_miss_vec_2 = 1'b0;
      end
    end else begin
      BTB_btb_is_miss_vec_2 = 1'b0;
    end
  end

  assign when_Predictor_l113_3 = (train_valid && train_taken);
  assign when_Predictor_l114_3 = ((BTB_source_pc_3 == train_pc) && BTB_valid[3]);
  always @(*) begin
    if(when_Predictor_l113_3) begin
      if(when_Predictor_l114_3) begin
        BTB_btb_is_hit_vec_3 = 1'b1;
      end else begin
        BTB_btb_is_hit_vec_3 = 1'b0;
      end
    end else begin
      BTB_btb_is_hit_vec_3 = 1'b0;
    end
  end

  assign when_Predictor_l119_3 = ((BTB_source_pc_3 != train_pc) || (! BTB_valid[3]));
  always @(*) begin
    if(when_Predictor_l113_3) begin
      if(when_Predictor_l119_3) begin
        BTB_btb_is_miss_vec_3 = 1'b1;
      end else begin
        BTB_btb_is_miss_vec_3 = 1'b0;
      end
    end else begin
      BTB_btb_is_miss_vec_3 = 1'b0;
    end
  end

  assign _zz_BTB_btb_write_index = (BTB_btb_is_hit_vec_1 || BTB_btb_is_hit_vec_3);
  assign _zz_BTB_btb_write_index_1 = (BTB_btb_is_hit_vec_2 || BTB_btb_is_hit_vec_3);
  assign BTB_btb_write_index = {_zz_BTB_btb_write_index_1,_zz_BTB_btb_write_index};
  assign _zz_130 = ({3'd0,1'b1} <<< BTB_btb_write_index);
  assign _zz_131 = ({3'd0,1'b1} <<< BTB_btb_write_index);
  assign _zz_132 = ({3'd0,1'b1} <<< BTB_btb_alloc_index_value);
  assign _zz_133 = ({3'd0,1'b1} <<< BTB_btb_alloc_index_value);
  assign RAS_ras_call_matched = (BTB_is_matched && BTB_is_call);
  assign RAS_ras_ret_matched = (BTB_is_matched && BTB_is_ret);
  assign when_Predictor_l169 = (train_valid && train_is_call);
  always @(*) begin
    if(when_Predictor_l169) begin
      RAS_ras_next_index_proven = (RAS_ras_curr_index_proven + 2'b01);
    end else begin
      if(when_Predictor_l172) begin
        RAS_ras_next_index_proven = (RAS_ras_curr_index_proven - 2'b01);
      end else begin
        RAS_ras_next_index_proven = RAS_ras_curr_index_proven;
      end
    end
  end

  assign when_Predictor_l172 = (train_valid && train_is_ret);
  assign when_Predictor_l180 = ((train_mispredicted && train_valid) && train_is_call);
  always @(*) begin
    if(when_Predictor_l180) begin
      RAS_ras_next_index = (RAS_ras_curr_index_proven + 2'b01);
    end else begin
      if(when_Predictor_l183) begin
        RAS_ras_next_index = (RAS_ras_curr_index_proven - 2'b01);
      end else begin
        if(RAS_ras_call_matched) begin
          RAS_ras_next_index = (RAS_ras_curr_index + 2'b01);
        end else begin
          if(RAS_ras_ret_matched) begin
            RAS_ras_next_index = (RAS_ras_curr_index - 2'b01);
          end else begin
            RAS_ras_next_index = RAS_ras_curr_index;
          end
        end
      end
    end
  end

  assign when_Predictor_l183 = ((train_mispredicted && train_valid) && train_is_ret);
  assign when_Predictor_l197 = ((train_mispredicted && train_valid) && train_is_call);
  assign _zz_134 = ({3'd0,1'b1} <<< RAS_ras_next_index);
  assign _zz_135 = _zz_134[0];
  assign _zz_136 = _zz_134[1];
  assign _zz_137 = _zz_134[2];
  assign _zz_138 = _zz_134[3];
  assign _zz_RAS_ras_regfile_0 = (train_pc + 64'h0000000000000004);
  assign _zz_RAS_ras_regfile_0_1 = (predict_pc + 64'h0000000000000004);
  assign when_Predictor_l205 = ((train_mispredicted && train_valid) && train_is_ret);
  assign RAS_ras_predict_pc = _zz_RAS_ras_predict_pc;
  assign predict_history = GSHARE_global_branch_history;
  assign predict_taken = (BTB_is_matched && (((GSHARE_pht_predict_taken || BTB_is_jmp) || BTB_is_call) || BTB_is_ret));
  assign predict_pc_next = (RAS_ras_ret_matched ? RAS_ras_predict_pc : ((BTB_is_matched && ((GSHARE_pht_predict_taken || BTB_is_jmp) || BTB_is_call)) ? BTB_target_pc_read : _zz_predict_pc_next));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      GSHARE_global_branch_history <= 7'h0;
      GSHARE_PHT_0 <= 2'b01;
      GSHARE_PHT_1 <= 2'b01;
      GSHARE_PHT_2 <= 2'b01;
      GSHARE_PHT_3 <= 2'b01;
      GSHARE_PHT_4 <= 2'b01;
      GSHARE_PHT_5 <= 2'b01;
      GSHARE_PHT_6 <= 2'b01;
      GSHARE_PHT_7 <= 2'b01;
      GSHARE_PHT_8 <= 2'b01;
      GSHARE_PHT_9 <= 2'b01;
      GSHARE_PHT_10 <= 2'b01;
      GSHARE_PHT_11 <= 2'b01;
      GSHARE_PHT_12 <= 2'b01;
      GSHARE_PHT_13 <= 2'b01;
      GSHARE_PHT_14 <= 2'b01;
      GSHARE_PHT_15 <= 2'b01;
      GSHARE_PHT_16 <= 2'b01;
      GSHARE_PHT_17 <= 2'b01;
      GSHARE_PHT_18 <= 2'b01;
      GSHARE_PHT_19 <= 2'b01;
      GSHARE_PHT_20 <= 2'b01;
      GSHARE_PHT_21 <= 2'b01;
      GSHARE_PHT_22 <= 2'b01;
      GSHARE_PHT_23 <= 2'b01;
      GSHARE_PHT_24 <= 2'b01;
      GSHARE_PHT_25 <= 2'b01;
      GSHARE_PHT_26 <= 2'b01;
      GSHARE_PHT_27 <= 2'b01;
      GSHARE_PHT_28 <= 2'b01;
      GSHARE_PHT_29 <= 2'b01;
      GSHARE_PHT_30 <= 2'b01;
      GSHARE_PHT_31 <= 2'b01;
      GSHARE_PHT_32 <= 2'b01;
      GSHARE_PHT_33 <= 2'b01;
      GSHARE_PHT_34 <= 2'b01;
      GSHARE_PHT_35 <= 2'b01;
      GSHARE_PHT_36 <= 2'b01;
      GSHARE_PHT_37 <= 2'b01;
      GSHARE_PHT_38 <= 2'b01;
      GSHARE_PHT_39 <= 2'b01;
      GSHARE_PHT_40 <= 2'b01;
      GSHARE_PHT_41 <= 2'b01;
      GSHARE_PHT_42 <= 2'b01;
      GSHARE_PHT_43 <= 2'b01;
      GSHARE_PHT_44 <= 2'b01;
      GSHARE_PHT_45 <= 2'b01;
      GSHARE_PHT_46 <= 2'b01;
      GSHARE_PHT_47 <= 2'b01;
      GSHARE_PHT_48 <= 2'b01;
      GSHARE_PHT_49 <= 2'b01;
      GSHARE_PHT_50 <= 2'b01;
      GSHARE_PHT_51 <= 2'b01;
      GSHARE_PHT_52 <= 2'b01;
      GSHARE_PHT_53 <= 2'b01;
      GSHARE_PHT_54 <= 2'b01;
      GSHARE_PHT_55 <= 2'b01;
      GSHARE_PHT_56 <= 2'b01;
      GSHARE_PHT_57 <= 2'b01;
      GSHARE_PHT_58 <= 2'b01;
      GSHARE_PHT_59 <= 2'b01;
      GSHARE_PHT_60 <= 2'b01;
      GSHARE_PHT_61 <= 2'b01;
      GSHARE_PHT_62 <= 2'b01;
      GSHARE_PHT_63 <= 2'b01;
      GSHARE_PHT_64 <= 2'b01;
      GSHARE_PHT_65 <= 2'b01;
      GSHARE_PHT_66 <= 2'b01;
      GSHARE_PHT_67 <= 2'b01;
      GSHARE_PHT_68 <= 2'b01;
      GSHARE_PHT_69 <= 2'b01;
      GSHARE_PHT_70 <= 2'b01;
      GSHARE_PHT_71 <= 2'b01;
      GSHARE_PHT_72 <= 2'b01;
      GSHARE_PHT_73 <= 2'b01;
      GSHARE_PHT_74 <= 2'b01;
      GSHARE_PHT_75 <= 2'b01;
      GSHARE_PHT_76 <= 2'b01;
      GSHARE_PHT_77 <= 2'b01;
      GSHARE_PHT_78 <= 2'b01;
      GSHARE_PHT_79 <= 2'b01;
      GSHARE_PHT_80 <= 2'b01;
      GSHARE_PHT_81 <= 2'b01;
      GSHARE_PHT_82 <= 2'b01;
      GSHARE_PHT_83 <= 2'b01;
      GSHARE_PHT_84 <= 2'b01;
      GSHARE_PHT_85 <= 2'b01;
      GSHARE_PHT_86 <= 2'b01;
      GSHARE_PHT_87 <= 2'b01;
      GSHARE_PHT_88 <= 2'b01;
      GSHARE_PHT_89 <= 2'b01;
      GSHARE_PHT_90 <= 2'b01;
      GSHARE_PHT_91 <= 2'b01;
      GSHARE_PHT_92 <= 2'b01;
      GSHARE_PHT_93 <= 2'b01;
      GSHARE_PHT_94 <= 2'b01;
      GSHARE_PHT_95 <= 2'b01;
      GSHARE_PHT_96 <= 2'b01;
      GSHARE_PHT_97 <= 2'b01;
      GSHARE_PHT_98 <= 2'b01;
      GSHARE_PHT_99 <= 2'b01;
      GSHARE_PHT_100 <= 2'b01;
      GSHARE_PHT_101 <= 2'b01;
      GSHARE_PHT_102 <= 2'b01;
      GSHARE_PHT_103 <= 2'b01;
      GSHARE_PHT_104 <= 2'b01;
      GSHARE_PHT_105 <= 2'b01;
      GSHARE_PHT_106 <= 2'b01;
      GSHARE_PHT_107 <= 2'b01;
      GSHARE_PHT_108 <= 2'b01;
      GSHARE_PHT_109 <= 2'b01;
      GSHARE_PHT_110 <= 2'b01;
      GSHARE_PHT_111 <= 2'b01;
      GSHARE_PHT_112 <= 2'b01;
      GSHARE_PHT_113 <= 2'b01;
      GSHARE_PHT_114 <= 2'b01;
      GSHARE_PHT_115 <= 2'b01;
      GSHARE_PHT_116 <= 2'b01;
      GSHARE_PHT_117 <= 2'b01;
      GSHARE_PHT_118 <= 2'b01;
      GSHARE_PHT_119 <= 2'b01;
      GSHARE_PHT_120 <= 2'b01;
      GSHARE_PHT_121 <= 2'b01;
      GSHARE_PHT_122 <= 2'b01;
      GSHARE_PHT_123 <= 2'b01;
      GSHARE_PHT_124 <= 2'b01;
      GSHARE_PHT_125 <= 2'b01;
      GSHARE_PHT_126 <= 2'b01;
      GSHARE_PHT_127 <= 2'b01;
      BTB_valid <= 4'b0000;
      BTB_source_pc_0 <= 64'h0;
      BTB_source_pc_1 <= 64'h0;
      BTB_source_pc_2 <= 64'h0;
      BTB_source_pc_3 <= 64'h0;
      BTB_call <= 4'b0000;
      BTB_ret <= 4'b0000;
      BTB_jmp <= 4'b0000;
      BTB_target_pc_0 <= 64'h0;
      BTB_target_pc_1 <= 64'h0;
      BTB_target_pc_2 <= 64'h0;
      BTB_target_pc_3 <= 64'h0;
      BTB_btb_alloc_index_value <= 2'b00;
      RAS_ras_curr_index <= 2'b00;
      RAS_ras_curr_index_proven <= 2'b00;
    end else begin
      if(train_valid) begin
        case(switch_Predictor_l38)
          2'b00 : begin
            if(train_taken) begin
              if(_zz_2) begin
                GSHARE_PHT_0 <= 2'b01;
              end
              if(_zz_3) begin
                GSHARE_PHT_1 <= 2'b01;
              end
              if(_zz_4) begin
                GSHARE_PHT_2 <= 2'b01;
              end
              if(_zz_5) begin
                GSHARE_PHT_3 <= 2'b01;
              end
              if(_zz_6) begin
                GSHARE_PHT_4 <= 2'b01;
              end
              if(_zz_7) begin
                GSHARE_PHT_5 <= 2'b01;
              end
              if(_zz_8) begin
                GSHARE_PHT_6 <= 2'b01;
              end
              if(_zz_9) begin
                GSHARE_PHT_7 <= 2'b01;
              end
              if(_zz_10) begin
                GSHARE_PHT_8 <= 2'b01;
              end
              if(_zz_11) begin
                GSHARE_PHT_9 <= 2'b01;
              end
              if(_zz_12) begin
                GSHARE_PHT_10 <= 2'b01;
              end
              if(_zz_13) begin
                GSHARE_PHT_11 <= 2'b01;
              end
              if(_zz_14) begin
                GSHARE_PHT_12 <= 2'b01;
              end
              if(_zz_15) begin
                GSHARE_PHT_13 <= 2'b01;
              end
              if(_zz_16) begin
                GSHARE_PHT_14 <= 2'b01;
              end
              if(_zz_17) begin
                GSHARE_PHT_15 <= 2'b01;
              end
              if(_zz_18) begin
                GSHARE_PHT_16 <= 2'b01;
              end
              if(_zz_19) begin
                GSHARE_PHT_17 <= 2'b01;
              end
              if(_zz_20) begin
                GSHARE_PHT_18 <= 2'b01;
              end
              if(_zz_21) begin
                GSHARE_PHT_19 <= 2'b01;
              end
              if(_zz_22) begin
                GSHARE_PHT_20 <= 2'b01;
              end
              if(_zz_23) begin
                GSHARE_PHT_21 <= 2'b01;
              end
              if(_zz_24) begin
                GSHARE_PHT_22 <= 2'b01;
              end
              if(_zz_25) begin
                GSHARE_PHT_23 <= 2'b01;
              end
              if(_zz_26) begin
                GSHARE_PHT_24 <= 2'b01;
              end
              if(_zz_27) begin
                GSHARE_PHT_25 <= 2'b01;
              end
              if(_zz_28) begin
                GSHARE_PHT_26 <= 2'b01;
              end
              if(_zz_29) begin
                GSHARE_PHT_27 <= 2'b01;
              end
              if(_zz_30) begin
                GSHARE_PHT_28 <= 2'b01;
              end
              if(_zz_31) begin
                GSHARE_PHT_29 <= 2'b01;
              end
              if(_zz_32) begin
                GSHARE_PHT_30 <= 2'b01;
              end
              if(_zz_33) begin
                GSHARE_PHT_31 <= 2'b01;
              end
              if(_zz_34) begin
                GSHARE_PHT_32 <= 2'b01;
              end
              if(_zz_35) begin
                GSHARE_PHT_33 <= 2'b01;
              end
              if(_zz_36) begin
                GSHARE_PHT_34 <= 2'b01;
              end
              if(_zz_37) begin
                GSHARE_PHT_35 <= 2'b01;
              end
              if(_zz_38) begin
                GSHARE_PHT_36 <= 2'b01;
              end
              if(_zz_39) begin
                GSHARE_PHT_37 <= 2'b01;
              end
              if(_zz_40) begin
                GSHARE_PHT_38 <= 2'b01;
              end
              if(_zz_41) begin
                GSHARE_PHT_39 <= 2'b01;
              end
              if(_zz_42) begin
                GSHARE_PHT_40 <= 2'b01;
              end
              if(_zz_43) begin
                GSHARE_PHT_41 <= 2'b01;
              end
              if(_zz_44) begin
                GSHARE_PHT_42 <= 2'b01;
              end
              if(_zz_45) begin
                GSHARE_PHT_43 <= 2'b01;
              end
              if(_zz_46) begin
                GSHARE_PHT_44 <= 2'b01;
              end
              if(_zz_47) begin
                GSHARE_PHT_45 <= 2'b01;
              end
              if(_zz_48) begin
                GSHARE_PHT_46 <= 2'b01;
              end
              if(_zz_49) begin
                GSHARE_PHT_47 <= 2'b01;
              end
              if(_zz_50) begin
                GSHARE_PHT_48 <= 2'b01;
              end
              if(_zz_51) begin
                GSHARE_PHT_49 <= 2'b01;
              end
              if(_zz_52) begin
                GSHARE_PHT_50 <= 2'b01;
              end
              if(_zz_53) begin
                GSHARE_PHT_51 <= 2'b01;
              end
              if(_zz_54) begin
                GSHARE_PHT_52 <= 2'b01;
              end
              if(_zz_55) begin
                GSHARE_PHT_53 <= 2'b01;
              end
              if(_zz_56) begin
                GSHARE_PHT_54 <= 2'b01;
              end
              if(_zz_57) begin
                GSHARE_PHT_55 <= 2'b01;
              end
              if(_zz_58) begin
                GSHARE_PHT_56 <= 2'b01;
              end
              if(_zz_59) begin
                GSHARE_PHT_57 <= 2'b01;
              end
              if(_zz_60) begin
                GSHARE_PHT_58 <= 2'b01;
              end
              if(_zz_61) begin
                GSHARE_PHT_59 <= 2'b01;
              end
              if(_zz_62) begin
                GSHARE_PHT_60 <= 2'b01;
              end
              if(_zz_63) begin
                GSHARE_PHT_61 <= 2'b01;
              end
              if(_zz_64) begin
                GSHARE_PHT_62 <= 2'b01;
              end
              if(_zz_65) begin
                GSHARE_PHT_63 <= 2'b01;
              end
              if(_zz_66) begin
                GSHARE_PHT_64 <= 2'b01;
              end
              if(_zz_67) begin
                GSHARE_PHT_65 <= 2'b01;
              end
              if(_zz_68) begin
                GSHARE_PHT_66 <= 2'b01;
              end
              if(_zz_69) begin
                GSHARE_PHT_67 <= 2'b01;
              end
              if(_zz_70) begin
                GSHARE_PHT_68 <= 2'b01;
              end
              if(_zz_71) begin
                GSHARE_PHT_69 <= 2'b01;
              end
              if(_zz_72) begin
                GSHARE_PHT_70 <= 2'b01;
              end
              if(_zz_73) begin
                GSHARE_PHT_71 <= 2'b01;
              end
              if(_zz_74) begin
                GSHARE_PHT_72 <= 2'b01;
              end
              if(_zz_75) begin
                GSHARE_PHT_73 <= 2'b01;
              end
              if(_zz_76) begin
                GSHARE_PHT_74 <= 2'b01;
              end
              if(_zz_77) begin
                GSHARE_PHT_75 <= 2'b01;
              end
              if(_zz_78) begin
                GSHARE_PHT_76 <= 2'b01;
              end
              if(_zz_79) begin
                GSHARE_PHT_77 <= 2'b01;
              end
              if(_zz_80) begin
                GSHARE_PHT_78 <= 2'b01;
              end
              if(_zz_81) begin
                GSHARE_PHT_79 <= 2'b01;
              end
              if(_zz_82) begin
                GSHARE_PHT_80 <= 2'b01;
              end
              if(_zz_83) begin
                GSHARE_PHT_81 <= 2'b01;
              end
              if(_zz_84) begin
                GSHARE_PHT_82 <= 2'b01;
              end
              if(_zz_85) begin
                GSHARE_PHT_83 <= 2'b01;
              end
              if(_zz_86) begin
                GSHARE_PHT_84 <= 2'b01;
              end
              if(_zz_87) begin
                GSHARE_PHT_85 <= 2'b01;
              end
              if(_zz_88) begin
                GSHARE_PHT_86 <= 2'b01;
              end
              if(_zz_89) begin
                GSHARE_PHT_87 <= 2'b01;
              end
              if(_zz_90) begin
                GSHARE_PHT_88 <= 2'b01;
              end
              if(_zz_91) begin
                GSHARE_PHT_89 <= 2'b01;
              end
              if(_zz_92) begin
                GSHARE_PHT_90 <= 2'b01;
              end
              if(_zz_93) begin
                GSHARE_PHT_91 <= 2'b01;
              end
              if(_zz_94) begin
                GSHARE_PHT_92 <= 2'b01;
              end
              if(_zz_95) begin
                GSHARE_PHT_93 <= 2'b01;
              end
              if(_zz_96) begin
                GSHARE_PHT_94 <= 2'b01;
              end
              if(_zz_97) begin
                GSHARE_PHT_95 <= 2'b01;
              end
              if(_zz_98) begin
                GSHARE_PHT_96 <= 2'b01;
              end
              if(_zz_99) begin
                GSHARE_PHT_97 <= 2'b01;
              end
              if(_zz_100) begin
                GSHARE_PHT_98 <= 2'b01;
              end
              if(_zz_101) begin
                GSHARE_PHT_99 <= 2'b01;
              end
              if(_zz_102) begin
                GSHARE_PHT_100 <= 2'b01;
              end
              if(_zz_103) begin
                GSHARE_PHT_101 <= 2'b01;
              end
              if(_zz_104) begin
                GSHARE_PHT_102 <= 2'b01;
              end
              if(_zz_105) begin
                GSHARE_PHT_103 <= 2'b01;
              end
              if(_zz_106) begin
                GSHARE_PHT_104 <= 2'b01;
              end
              if(_zz_107) begin
                GSHARE_PHT_105 <= 2'b01;
              end
              if(_zz_108) begin
                GSHARE_PHT_106 <= 2'b01;
              end
              if(_zz_109) begin
                GSHARE_PHT_107 <= 2'b01;
              end
              if(_zz_110) begin
                GSHARE_PHT_108 <= 2'b01;
              end
              if(_zz_111) begin
                GSHARE_PHT_109 <= 2'b01;
              end
              if(_zz_112) begin
                GSHARE_PHT_110 <= 2'b01;
              end
              if(_zz_113) begin
                GSHARE_PHT_111 <= 2'b01;
              end
              if(_zz_114) begin
                GSHARE_PHT_112 <= 2'b01;
              end
              if(_zz_115) begin
                GSHARE_PHT_113 <= 2'b01;
              end
              if(_zz_116) begin
                GSHARE_PHT_114 <= 2'b01;
              end
              if(_zz_117) begin
                GSHARE_PHT_115 <= 2'b01;
              end
              if(_zz_118) begin
                GSHARE_PHT_116 <= 2'b01;
              end
              if(_zz_119) begin
                GSHARE_PHT_117 <= 2'b01;
              end
              if(_zz_120) begin
                GSHARE_PHT_118 <= 2'b01;
              end
              if(_zz_121) begin
                GSHARE_PHT_119 <= 2'b01;
              end
              if(_zz_122) begin
                GSHARE_PHT_120 <= 2'b01;
              end
              if(_zz_123) begin
                GSHARE_PHT_121 <= 2'b01;
              end
              if(_zz_124) begin
                GSHARE_PHT_122 <= 2'b01;
              end
              if(_zz_125) begin
                GSHARE_PHT_123 <= 2'b01;
              end
              if(_zz_126) begin
                GSHARE_PHT_124 <= 2'b01;
              end
              if(_zz_127) begin
                GSHARE_PHT_125 <= 2'b01;
              end
              if(_zz_128) begin
                GSHARE_PHT_126 <= 2'b01;
              end
              if(_zz_129) begin
                GSHARE_PHT_127 <= 2'b01;
              end
            end else begin
              if(_zz_2) begin
                GSHARE_PHT_0 <= 2'b00;
              end
              if(_zz_3) begin
                GSHARE_PHT_1 <= 2'b00;
              end
              if(_zz_4) begin
                GSHARE_PHT_2 <= 2'b00;
              end
              if(_zz_5) begin
                GSHARE_PHT_3 <= 2'b00;
              end
              if(_zz_6) begin
                GSHARE_PHT_4 <= 2'b00;
              end
              if(_zz_7) begin
                GSHARE_PHT_5 <= 2'b00;
              end
              if(_zz_8) begin
                GSHARE_PHT_6 <= 2'b00;
              end
              if(_zz_9) begin
                GSHARE_PHT_7 <= 2'b00;
              end
              if(_zz_10) begin
                GSHARE_PHT_8 <= 2'b00;
              end
              if(_zz_11) begin
                GSHARE_PHT_9 <= 2'b00;
              end
              if(_zz_12) begin
                GSHARE_PHT_10 <= 2'b00;
              end
              if(_zz_13) begin
                GSHARE_PHT_11 <= 2'b00;
              end
              if(_zz_14) begin
                GSHARE_PHT_12 <= 2'b00;
              end
              if(_zz_15) begin
                GSHARE_PHT_13 <= 2'b00;
              end
              if(_zz_16) begin
                GSHARE_PHT_14 <= 2'b00;
              end
              if(_zz_17) begin
                GSHARE_PHT_15 <= 2'b00;
              end
              if(_zz_18) begin
                GSHARE_PHT_16 <= 2'b00;
              end
              if(_zz_19) begin
                GSHARE_PHT_17 <= 2'b00;
              end
              if(_zz_20) begin
                GSHARE_PHT_18 <= 2'b00;
              end
              if(_zz_21) begin
                GSHARE_PHT_19 <= 2'b00;
              end
              if(_zz_22) begin
                GSHARE_PHT_20 <= 2'b00;
              end
              if(_zz_23) begin
                GSHARE_PHT_21 <= 2'b00;
              end
              if(_zz_24) begin
                GSHARE_PHT_22 <= 2'b00;
              end
              if(_zz_25) begin
                GSHARE_PHT_23 <= 2'b00;
              end
              if(_zz_26) begin
                GSHARE_PHT_24 <= 2'b00;
              end
              if(_zz_27) begin
                GSHARE_PHT_25 <= 2'b00;
              end
              if(_zz_28) begin
                GSHARE_PHT_26 <= 2'b00;
              end
              if(_zz_29) begin
                GSHARE_PHT_27 <= 2'b00;
              end
              if(_zz_30) begin
                GSHARE_PHT_28 <= 2'b00;
              end
              if(_zz_31) begin
                GSHARE_PHT_29 <= 2'b00;
              end
              if(_zz_32) begin
                GSHARE_PHT_30 <= 2'b00;
              end
              if(_zz_33) begin
                GSHARE_PHT_31 <= 2'b00;
              end
              if(_zz_34) begin
                GSHARE_PHT_32 <= 2'b00;
              end
              if(_zz_35) begin
                GSHARE_PHT_33 <= 2'b00;
              end
              if(_zz_36) begin
                GSHARE_PHT_34 <= 2'b00;
              end
              if(_zz_37) begin
                GSHARE_PHT_35 <= 2'b00;
              end
              if(_zz_38) begin
                GSHARE_PHT_36 <= 2'b00;
              end
              if(_zz_39) begin
                GSHARE_PHT_37 <= 2'b00;
              end
              if(_zz_40) begin
                GSHARE_PHT_38 <= 2'b00;
              end
              if(_zz_41) begin
                GSHARE_PHT_39 <= 2'b00;
              end
              if(_zz_42) begin
                GSHARE_PHT_40 <= 2'b00;
              end
              if(_zz_43) begin
                GSHARE_PHT_41 <= 2'b00;
              end
              if(_zz_44) begin
                GSHARE_PHT_42 <= 2'b00;
              end
              if(_zz_45) begin
                GSHARE_PHT_43 <= 2'b00;
              end
              if(_zz_46) begin
                GSHARE_PHT_44 <= 2'b00;
              end
              if(_zz_47) begin
                GSHARE_PHT_45 <= 2'b00;
              end
              if(_zz_48) begin
                GSHARE_PHT_46 <= 2'b00;
              end
              if(_zz_49) begin
                GSHARE_PHT_47 <= 2'b00;
              end
              if(_zz_50) begin
                GSHARE_PHT_48 <= 2'b00;
              end
              if(_zz_51) begin
                GSHARE_PHT_49 <= 2'b00;
              end
              if(_zz_52) begin
                GSHARE_PHT_50 <= 2'b00;
              end
              if(_zz_53) begin
                GSHARE_PHT_51 <= 2'b00;
              end
              if(_zz_54) begin
                GSHARE_PHT_52 <= 2'b00;
              end
              if(_zz_55) begin
                GSHARE_PHT_53 <= 2'b00;
              end
              if(_zz_56) begin
                GSHARE_PHT_54 <= 2'b00;
              end
              if(_zz_57) begin
                GSHARE_PHT_55 <= 2'b00;
              end
              if(_zz_58) begin
                GSHARE_PHT_56 <= 2'b00;
              end
              if(_zz_59) begin
                GSHARE_PHT_57 <= 2'b00;
              end
              if(_zz_60) begin
                GSHARE_PHT_58 <= 2'b00;
              end
              if(_zz_61) begin
                GSHARE_PHT_59 <= 2'b00;
              end
              if(_zz_62) begin
                GSHARE_PHT_60 <= 2'b00;
              end
              if(_zz_63) begin
                GSHARE_PHT_61 <= 2'b00;
              end
              if(_zz_64) begin
                GSHARE_PHT_62 <= 2'b00;
              end
              if(_zz_65) begin
                GSHARE_PHT_63 <= 2'b00;
              end
              if(_zz_66) begin
                GSHARE_PHT_64 <= 2'b00;
              end
              if(_zz_67) begin
                GSHARE_PHT_65 <= 2'b00;
              end
              if(_zz_68) begin
                GSHARE_PHT_66 <= 2'b00;
              end
              if(_zz_69) begin
                GSHARE_PHT_67 <= 2'b00;
              end
              if(_zz_70) begin
                GSHARE_PHT_68 <= 2'b00;
              end
              if(_zz_71) begin
                GSHARE_PHT_69 <= 2'b00;
              end
              if(_zz_72) begin
                GSHARE_PHT_70 <= 2'b00;
              end
              if(_zz_73) begin
                GSHARE_PHT_71 <= 2'b00;
              end
              if(_zz_74) begin
                GSHARE_PHT_72 <= 2'b00;
              end
              if(_zz_75) begin
                GSHARE_PHT_73 <= 2'b00;
              end
              if(_zz_76) begin
                GSHARE_PHT_74 <= 2'b00;
              end
              if(_zz_77) begin
                GSHARE_PHT_75 <= 2'b00;
              end
              if(_zz_78) begin
                GSHARE_PHT_76 <= 2'b00;
              end
              if(_zz_79) begin
                GSHARE_PHT_77 <= 2'b00;
              end
              if(_zz_80) begin
                GSHARE_PHT_78 <= 2'b00;
              end
              if(_zz_81) begin
                GSHARE_PHT_79 <= 2'b00;
              end
              if(_zz_82) begin
                GSHARE_PHT_80 <= 2'b00;
              end
              if(_zz_83) begin
                GSHARE_PHT_81 <= 2'b00;
              end
              if(_zz_84) begin
                GSHARE_PHT_82 <= 2'b00;
              end
              if(_zz_85) begin
                GSHARE_PHT_83 <= 2'b00;
              end
              if(_zz_86) begin
                GSHARE_PHT_84 <= 2'b00;
              end
              if(_zz_87) begin
                GSHARE_PHT_85 <= 2'b00;
              end
              if(_zz_88) begin
                GSHARE_PHT_86 <= 2'b00;
              end
              if(_zz_89) begin
                GSHARE_PHT_87 <= 2'b00;
              end
              if(_zz_90) begin
                GSHARE_PHT_88 <= 2'b00;
              end
              if(_zz_91) begin
                GSHARE_PHT_89 <= 2'b00;
              end
              if(_zz_92) begin
                GSHARE_PHT_90 <= 2'b00;
              end
              if(_zz_93) begin
                GSHARE_PHT_91 <= 2'b00;
              end
              if(_zz_94) begin
                GSHARE_PHT_92 <= 2'b00;
              end
              if(_zz_95) begin
                GSHARE_PHT_93 <= 2'b00;
              end
              if(_zz_96) begin
                GSHARE_PHT_94 <= 2'b00;
              end
              if(_zz_97) begin
                GSHARE_PHT_95 <= 2'b00;
              end
              if(_zz_98) begin
                GSHARE_PHT_96 <= 2'b00;
              end
              if(_zz_99) begin
                GSHARE_PHT_97 <= 2'b00;
              end
              if(_zz_100) begin
                GSHARE_PHT_98 <= 2'b00;
              end
              if(_zz_101) begin
                GSHARE_PHT_99 <= 2'b00;
              end
              if(_zz_102) begin
                GSHARE_PHT_100 <= 2'b00;
              end
              if(_zz_103) begin
                GSHARE_PHT_101 <= 2'b00;
              end
              if(_zz_104) begin
                GSHARE_PHT_102 <= 2'b00;
              end
              if(_zz_105) begin
                GSHARE_PHT_103 <= 2'b00;
              end
              if(_zz_106) begin
                GSHARE_PHT_104 <= 2'b00;
              end
              if(_zz_107) begin
                GSHARE_PHT_105 <= 2'b00;
              end
              if(_zz_108) begin
                GSHARE_PHT_106 <= 2'b00;
              end
              if(_zz_109) begin
                GSHARE_PHT_107 <= 2'b00;
              end
              if(_zz_110) begin
                GSHARE_PHT_108 <= 2'b00;
              end
              if(_zz_111) begin
                GSHARE_PHT_109 <= 2'b00;
              end
              if(_zz_112) begin
                GSHARE_PHT_110 <= 2'b00;
              end
              if(_zz_113) begin
                GSHARE_PHT_111 <= 2'b00;
              end
              if(_zz_114) begin
                GSHARE_PHT_112 <= 2'b00;
              end
              if(_zz_115) begin
                GSHARE_PHT_113 <= 2'b00;
              end
              if(_zz_116) begin
                GSHARE_PHT_114 <= 2'b00;
              end
              if(_zz_117) begin
                GSHARE_PHT_115 <= 2'b00;
              end
              if(_zz_118) begin
                GSHARE_PHT_116 <= 2'b00;
              end
              if(_zz_119) begin
                GSHARE_PHT_117 <= 2'b00;
              end
              if(_zz_120) begin
                GSHARE_PHT_118 <= 2'b00;
              end
              if(_zz_121) begin
                GSHARE_PHT_119 <= 2'b00;
              end
              if(_zz_122) begin
                GSHARE_PHT_120 <= 2'b00;
              end
              if(_zz_123) begin
                GSHARE_PHT_121 <= 2'b00;
              end
              if(_zz_124) begin
                GSHARE_PHT_122 <= 2'b00;
              end
              if(_zz_125) begin
                GSHARE_PHT_123 <= 2'b00;
              end
              if(_zz_126) begin
                GSHARE_PHT_124 <= 2'b00;
              end
              if(_zz_127) begin
                GSHARE_PHT_125 <= 2'b00;
              end
              if(_zz_128) begin
                GSHARE_PHT_126 <= 2'b00;
              end
              if(_zz_129) begin
                GSHARE_PHT_127 <= 2'b00;
              end
            end
          end
          2'b01 : begin
            if(train_taken) begin
              if(_zz_2) begin
                GSHARE_PHT_0 <= 2'b10;
              end
              if(_zz_3) begin
                GSHARE_PHT_1 <= 2'b10;
              end
              if(_zz_4) begin
                GSHARE_PHT_2 <= 2'b10;
              end
              if(_zz_5) begin
                GSHARE_PHT_3 <= 2'b10;
              end
              if(_zz_6) begin
                GSHARE_PHT_4 <= 2'b10;
              end
              if(_zz_7) begin
                GSHARE_PHT_5 <= 2'b10;
              end
              if(_zz_8) begin
                GSHARE_PHT_6 <= 2'b10;
              end
              if(_zz_9) begin
                GSHARE_PHT_7 <= 2'b10;
              end
              if(_zz_10) begin
                GSHARE_PHT_8 <= 2'b10;
              end
              if(_zz_11) begin
                GSHARE_PHT_9 <= 2'b10;
              end
              if(_zz_12) begin
                GSHARE_PHT_10 <= 2'b10;
              end
              if(_zz_13) begin
                GSHARE_PHT_11 <= 2'b10;
              end
              if(_zz_14) begin
                GSHARE_PHT_12 <= 2'b10;
              end
              if(_zz_15) begin
                GSHARE_PHT_13 <= 2'b10;
              end
              if(_zz_16) begin
                GSHARE_PHT_14 <= 2'b10;
              end
              if(_zz_17) begin
                GSHARE_PHT_15 <= 2'b10;
              end
              if(_zz_18) begin
                GSHARE_PHT_16 <= 2'b10;
              end
              if(_zz_19) begin
                GSHARE_PHT_17 <= 2'b10;
              end
              if(_zz_20) begin
                GSHARE_PHT_18 <= 2'b10;
              end
              if(_zz_21) begin
                GSHARE_PHT_19 <= 2'b10;
              end
              if(_zz_22) begin
                GSHARE_PHT_20 <= 2'b10;
              end
              if(_zz_23) begin
                GSHARE_PHT_21 <= 2'b10;
              end
              if(_zz_24) begin
                GSHARE_PHT_22 <= 2'b10;
              end
              if(_zz_25) begin
                GSHARE_PHT_23 <= 2'b10;
              end
              if(_zz_26) begin
                GSHARE_PHT_24 <= 2'b10;
              end
              if(_zz_27) begin
                GSHARE_PHT_25 <= 2'b10;
              end
              if(_zz_28) begin
                GSHARE_PHT_26 <= 2'b10;
              end
              if(_zz_29) begin
                GSHARE_PHT_27 <= 2'b10;
              end
              if(_zz_30) begin
                GSHARE_PHT_28 <= 2'b10;
              end
              if(_zz_31) begin
                GSHARE_PHT_29 <= 2'b10;
              end
              if(_zz_32) begin
                GSHARE_PHT_30 <= 2'b10;
              end
              if(_zz_33) begin
                GSHARE_PHT_31 <= 2'b10;
              end
              if(_zz_34) begin
                GSHARE_PHT_32 <= 2'b10;
              end
              if(_zz_35) begin
                GSHARE_PHT_33 <= 2'b10;
              end
              if(_zz_36) begin
                GSHARE_PHT_34 <= 2'b10;
              end
              if(_zz_37) begin
                GSHARE_PHT_35 <= 2'b10;
              end
              if(_zz_38) begin
                GSHARE_PHT_36 <= 2'b10;
              end
              if(_zz_39) begin
                GSHARE_PHT_37 <= 2'b10;
              end
              if(_zz_40) begin
                GSHARE_PHT_38 <= 2'b10;
              end
              if(_zz_41) begin
                GSHARE_PHT_39 <= 2'b10;
              end
              if(_zz_42) begin
                GSHARE_PHT_40 <= 2'b10;
              end
              if(_zz_43) begin
                GSHARE_PHT_41 <= 2'b10;
              end
              if(_zz_44) begin
                GSHARE_PHT_42 <= 2'b10;
              end
              if(_zz_45) begin
                GSHARE_PHT_43 <= 2'b10;
              end
              if(_zz_46) begin
                GSHARE_PHT_44 <= 2'b10;
              end
              if(_zz_47) begin
                GSHARE_PHT_45 <= 2'b10;
              end
              if(_zz_48) begin
                GSHARE_PHT_46 <= 2'b10;
              end
              if(_zz_49) begin
                GSHARE_PHT_47 <= 2'b10;
              end
              if(_zz_50) begin
                GSHARE_PHT_48 <= 2'b10;
              end
              if(_zz_51) begin
                GSHARE_PHT_49 <= 2'b10;
              end
              if(_zz_52) begin
                GSHARE_PHT_50 <= 2'b10;
              end
              if(_zz_53) begin
                GSHARE_PHT_51 <= 2'b10;
              end
              if(_zz_54) begin
                GSHARE_PHT_52 <= 2'b10;
              end
              if(_zz_55) begin
                GSHARE_PHT_53 <= 2'b10;
              end
              if(_zz_56) begin
                GSHARE_PHT_54 <= 2'b10;
              end
              if(_zz_57) begin
                GSHARE_PHT_55 <= 2'b10;
              end
              if(_zz_58) begin
                GSHARE_PHT_56 <= 2'b10;
              end
              if(_zz_59) begin
                GSHARE_PHT_57 <= 2'b10;
              end
              if(_zz_60) begin
                GSHARE_PHT_58 <= 2'b10;
              end
              if(_zz_61) begin
                GSHARE_PHT_59 <= 2'b10;
              end
              if(_zz_62) begin
                GSHARE_PHT_60 <= 2'b10;
              end
              if(_zz_63) begin
                GSHARE_PHT_61 <= 2'b10;
              end
              if(_zz_64) begin
                GSHARE_PHT_62 <= 2'b10;
              end
              if(_zz_65) begin
                GSHARE_PHT_63 <= 2'b10;
              end
              if(_zz_66) begin
                GSHARE_PHT_64 <= 2'b10;
              end
              if(_zz_67) begin
                GSHARE_PHT_65 <= 2'b10;
              end
              if(_zz_68) begin
                GSHARE_PHT_66 <= 2'b10;
              end
              if(_zz_69) begin
                GSHARE_PHT_67 <= 2'b10;
              end
              if(_zz_70) begin
                GSHARE_PHT_68 <= 2'b10;
              end
              if(_zz_71) begin
                GSHARE_PHT_69 <= 2'b10;
              end
              if(_zz_72) begin
                GSHARE_PHT_70 <= 2'b10;
              end
              if(_zz_73) begin
                GSHARE_PHT_71 <= 2'b10;
              end
              if(_zz_74) begin
                GSHARE_PHT_72 <= 2'b10;
              end
              if(_zz_75) begin
                GSHARE_PHT_73 <= 2'b10;
              end
              if(_zz_76) begin
                GSHARE_PHT_74 <= 2'b10;
              end
              if(_zz_77) begin
                GSHARE_PHT_75 <= 2'b10;
              end
              if(_zz_78) begin
                GSHARE_PHT_76 <= 2'b10;
              end
              if(_zz_79) begin
                GSHARE_PHT_77 <= 2'b10;
              end
              if(_zz_80) begin
                GSHARE_PHT_78 <= 2'b10;
              end
              if(_zz_81) begin
                GSHARE_PHT_79 <= 2'b10;
              end
              if(_zz_82) begin
                GSHARE_PHT_80 <= 2'b10;
              end
              if(_zz_83) begin
                GSHARE_PHT_81 <= 2'b10;
              end
              if(_zz_84) begin
                GSHARE_PHT_82 <= 2'b10;
              end
              if(_zz_85) begin
                GSHARE_PHT_83 <= 2'b10;
              end
              if(_zz_86) begin
                GSHARE_PHT_84 <= 2'b10;
              end
              if(_zz_87) begin
                GSHARE_PHT_85 <= 2'b10;
              end
              if(_zz_88) begin
                GSHARE_PHT_86 <= 2'b10;
              end
              if(_zz_89) begin
                GSHARE_PHT_87 <= 2'b10;
              end
              if(_zz_90) begin
                GSHARE_PHT_88 <= 2'b10;
              end
              if(_zz_91) begin
                GSHARE_PHT_89 <= 2'b10;
              end
              if(_zz_92) begin
                GSHARE_PHT_90 <= 2'b10;
              end
              if(_zz_93) begin
                GSHARE_PHT_91 <= 2'b10;
              end
              if(_zz_94) begin
                GSHARE_PHT_92 <= 2'b10;
              end
              if(_zz_95) begin
                GSHARE_PHT_93 <= 2'b10;
              end
              if(_zz_96) begin
                GSHARE_PHT_94 <= 2'b10;
              end
              if(_zz_97) begin
                GSHARE_PHT_95 <= 2'b10;
              end
              if(_zz_98) begin
                GSHARE_PHT_96 <= 2'b10;
              end
              if(_zz_99) begin
                GSHARE_PHT_97 <= 2'b10;
              end
              if(_zz_100) begin
                GSHARE_PHT_98 <= 2'b10;
              end
              if(_zz_101) begin
                GSHARE_PHT_99 <= 2'b10;
              end
              if(_zz_102) begin
                GSHARE_PHT_100 <= 2'b10;
              end
              if(_zz_103) begin
                GSHARE_PHT_101 <= 2'b10;
              end
              if(_zz_104) begin
                GSHARE_PHT_102 <= 2'b10;
              end
              if(_zz_105) begin
                GSHARE_PHT_103 <= 2'b10;
              end
              if(_zz_106) begin
                GSHARE_PHT_104 <= 2'b10;
              end
              if(_zz_107) begin
                GSHARE_PHT_105 <= 2'b10;
              end
              if(_zz_108) begin
                GSHARE_PHT_106 <= 2'b10;
              end
              if(_zz_109) begin
                GSHARE_PHT_107 <= 2'b10;
              end
              if(_zz_110) begin
                GSHARE_PHT_108 <= 2'b10;
              end
              if(_zz_111) begin
                GSHARE_PHT_109 <= 2'b10;
              end
              if(_zz_112) begin
                GSHARE_PHT_110 <= 2'b10;
              end
              if(_zz_113) begin
                GSHARE_PHT_111 <= 2'b10;
              end
              if(_zz_114) begin
                GSHARE_PHT_112 <= 2'b10;
              end
              if(_zz_115) begin
                GSHARE_PHT_113 <= 2'b10;
              end
              if(_zz_116) begin
                GSHARE_PHT_114 <= 2'b10;
              end
              if(_zz_117) begin
                GSHARE_PHT_115 <= 2'b10;
              end
              if(_zz_118) begin
                GSHARE_PHT_116 <= 2'b10;
              end
              if(_zz_119) begin
                GSHARE_PHT_117 <= 2'b10;
              end
              if(_zz_120) begin
                GSHARE_PHT_118 <= 2'b10;
              end
              if(_zz_121) begin
                GSHARE_PHT_119 <= 2'b10;
              end
              if(_zz_122) begin
                GSHARE_PHT_120 <= 2'b10;
              end
              if(_zz_123) begin
                GSHARE_PHT_121 <= 2'b10;
              end
              if(_zz_124) begin
                GSHARE_PHT_122 <= 2'b10;
              end
              if(_zz_125) begin
                GSHARE_PHT_123 <= 2'b10;
              end
              if(_zz_126) begin
                GSHARE_PHT_124 <= 2'b10;
              end
              if(_zz_127) begin
                GSHARE_PHT_125 <= 2'b10;
              end
              if(_zz_128) begin
                GSHARE_PHT_126 <= 2'b10;
              end
              if(_zz_129) begin
                GSHARE_PHT_127 <= 2'b10;
              end
            end else begin
              if(_zz_2) begin
                GSHARE_PHT_0 <= 2'b00;
              end
              if(_zz_3) begin
                GSHARE_PHT_1 <= 2'b00;
              end
              if(_zz_4) begin
                GSHARE_PHT_2 <= 2'b00;
              end
              if(_zz_5) begin
                GSHARE_PHT_3 <= 2'b00;
              end
              if(_zz_6) begin
                GSHARE_PHT_4 <= 2'b00;
              end
              if(_zz_7) begin
                GSHARE_PHT_5 <= 2'b00;
              end
              if(_zz_8) begin
                GSHARE_PHT_6 <= 2'b00;
              end
              if(_zz_9) begin
                GSHARE_PHT_7 <= 2'b00;
              end
              if(_zz_10) begin
                GSHARE_PHT_8 <= 2'b00;
              end
              if(_zz_11) begin
                GSHARE_PHT_9 <= 2'b00;
              end
              if(_zz_12) begin
                GSHARE_PHT_10 <= 2'b00;
              end
              if(_zz_13) begin
                GSHARE_PHT_11 <= 2'b00;
              end
              if(_zz_14) begin
                GSHARE_PHT_12 <= 2'b00;
              end
              if(_zz_15) begin
                GSHARE_PHT_13 <= 2'b00;
              end
              if(_zz_16) begin
                GSHARE_PHT_14 <= 2'b00;
              end
              if(_zz_17) begin
                GSHARE_PHT_15 <= 2'b00;
              end
              if(_zz_18) begin
                GSHARE_PHT_16 <= 2'b00;
              end
              if(_zz_19) begin
                GSHARE_PHT_17 <= 2'b00;
              end
              if(_zz_20) begin
                GSHARE_PHT_18 <= 2'b00;
              end
              if(_zz_21) begin
                GSHARE_PHT_19 <= 2'b00;
              end
              if(_zz_22) begin
                GSHARE_PHT_20 <= 2'b00;
              end
              if(_zz_23) begin
                GSHARE_PHT_21 <= 2'b00;
              end
              if(_zz_24) begin
                GSHARE_PHT_22 <= 2'b00;
              end
              if(_zz_25) begin
                GSHARE_PHT_23 <= 2'b00;
              end
              if(_zz_26) begin
                GSHARE_PHT_24 <= 2'b00;
              end
              if(_zz_27) begin
                GSHARE_PHT_25 <= 2'b00;
              end
              if(_zz_28) begin
                GSHARE_PHT_26 <= 2'b00;
              end
              if(_zz_29) begin
                GSHARE_PHT_27 <= 2'b00;
              end
              if(_zz_30) begin
                GSHARE_PHT_28 <= 2'b00;
              end
              if(_zz_31) begin
                GSHARE_PHT_29 <= 2'b00;
              end
              if(_zz_32) begin
                GSHARE_PHT_30 <= 2'b00;
              end
              if(_zz_33) begin
                GSHARE_PHT_31 <= 2'b00;
              end
              if(_zz_34) begin
                GSHARE_PHT_32 <= 2'b00;
              end
              if(_zz_35) begin
                GSHARE_PHT_33 <= 2'b00;
              end
              if(_zz_36) begin
                GSHARE_PHT_34 <= 2'b00;
              end
              if(_zz_37) begin
                GSHARE_PHT_35 <= 2'b00;
              end
              if(_zz_38) begin
                GSHARE_PHT_36 <= 2'b00;
              end
              if(_zz_39) begin
                GSHARE_PHT_37 <= 2'b00;
              end
              if(_zz_40) begin
                GSHARE_PHT_38 <= 2'b00;
              end
              if(_zz_41) begin
                GSHARE_PHT_39 <= 2'b00;
              end
              if(_zz_42) begin
                GSHARE_PHT_40 <= 2'b00;
              end
              if(_zz_43) begin
                GSHARE_PHT_41 <= 2'b00;
              end
              if(_zz_44) begin
                GSHARE_PHT_42 <= 2'b00;
              end
              if(_zz_45) begin
                GSHARE_PHT_43 <= 2'b00;
              end
              if(_zz_46) begin
                GSHARE_PHT_44 <= 2'b00;
              end
              if(_zz_47) begin
                GSHARE_PHT_45 <= 2'b00;
              end
              if(_zz_48) begin
                GSHARE_PHT_46 <= 2'b00;
              end
              if(_zz_49) begin
                GSHARE_PHT_47 <= 2'b00;
              end
              if(_zz_50) begin
                GSHARE_PHT_48 <= 2'b00;
              end
              if(_zz_51) begin
                GSHARE_PHT_49 <= 2'b00;
              end
              if(_zz_52) begin
                GSHARE_PHT_50 <= 2'b00;
              end
              if(_zz_53) begin
                GSHARE_PHT_51 <= 2'b00;
              end
              if(_zz_54) begin
                GSHARE_PHT_52 <= 2'b00;
              end
              if(_zz_55) begin
                GSHARE_PHT_53 <= 2'b00;
              end
              if(_zz_56) begin
                GSHARE_PHT_54 <= 2'b00;
              end
              if(_zz_57) begin
                GSHARE_PHT_55 <= 2'b00;
              end
              if(_zz_58) begin
                GSHARE_PHT_56 <= 2'b00;
              end
              if(_zz_59) begin
                GSHARE_PHT_57 <= 2'b00;
              end
              if(_zz_60) begin
                GSHARE_PHT_58 <= 2'b00;
              end
              if(_zz_61) begin
                GSHARE_PHT_59 <= 2'b00;
              end
              if(_zz_62) begin
                GSHARE_PHT_60 <= 2'b00;
              end
              if(_zz_63) begin
                GSHARE_PHT_61 <= 2'b00;
              end
              if(_zz_64) begin
                GSHARE_PHT_62 <= 2'b00;
              end
              if(_zz_65) begin
                GSHARE_PHT_63 <= 2'b00;
              end
              if(_zz_66) begin
                GSHARE_PHT_64 <= 2'b00;
              end
              if(_zz_67) begin
                GSHARE_PHT_65 <= 2'b00;
              end
              if(_zz_68) begin
                GSHARE_PHT_66 <= 2'b00;
              end
              if(_zz_69) begin
                GSHARE_PHT_67 <= 2'b00;
              end
              if(_zz_70) begin
                GSHARE_PHT_68 <= 2'b00;
              end
              if(_zz_71) begin
                GSHARE_PHT_69 <= 2'b00;
              end
              if(_zz_72) begin
                GSHARE_PHT_70 <= 2'b00;
              end
              if(_zz_73) begin
                GSHARE_PHT_71 <= 2'b00;
              end
              if(_zz_74) begin
                GSHARE_PHT_72 <= 2'b00;
              end
              if(_zz_75) begin
                GSHARE_PHT_73 <= 2'b00;
              end
              if(_zz_76) begin
                GSHARE_PHT_74 <= 2'b00;
              end
              if(_zz_77) begin
                GSHARE_PHT_75 <= 2'b00;
              end
              if(_zz_78) begin
                GSHARE_PHT_76 <= 2'b00;
              end
              if(_zz_79) begin
                GSHARE_PHT_77 <= 2'b00;
              end
              if(_zz_80) begin
                GSHARE_PHT_78 <= 2'b00;
              end
              if(_zz_81) begin
                GSHARE_PHT_79 <= 2'b00;
              end
              if(_zz_82) begin
                GSHARE_PHT_80 <= 2'b00;
              end
              if(_zz_83) begin
                GSHARE_PHT_81 <= 2'b00;
              end
              if(_zz_84) begin
                GSHARE_PHT_82 <= 2'b00;
              end
              if(_zz_85) begin
                GSHARE_PHT_83 <= 2'b00;
              end
              if(_zz_86) begin
                GSHARE_PHT_84 <= 2'b00;
              end
              if(_zz_87) begin
                GSHARE_PHT_85 <= 2'b00;
              end
              if(_zz_88) begin
                GSHARE_PHT_86 <= 2'b00;
              end
              if(_zz_89) begin
                GSHARE_PHT_87 <= 2'b00;
              end
              if(_zz_90) begin
                GSHARE_PHT_88 <= 2'b00;
              end
              if(_zz_91) begin
                GSHARE_PHT_89 <= 2'b00;
              end
              if(_zz_92) begin
                GSHARE_PHT_90 <= 2'b00;
              end
              if(_zz_93) begin
                GSHARE_PHT_91 <= 2'b00;
              end
              if(_zz_94) begin
                GSHARE_PHT_92 <= 2'b00;
              end
              if(_zz_95) begin
                GSHARE_PHT_93 <= 2'b00;
              end
              if(_zz_96) begin
                GSHARE_PHT_94 <= 2'b00;
              end
              if(_zz_97) begin
                GSHARE_PHT_95 <= 2'b00;
              end
              if(_zz_98) begin
                GSHARE_PHT_96 <= 2'b00;
              end
              if(_zz_99) begin
                GSHARE_PHT_97 <= 2'b00;
              end
              if(_zz_100) begin
                GSHARE_PHT_98 <= 2'b00;
              end
              if(_zz_101) begin
                GSHARE_PHT_99 <= 2'b00;
              end
              if(_zz_102) begin
                GSHARE_PHT_100 <= 2'b00;
              end
              if(_zz_103) begin
                GSHARE_PHT_101 <= 2'b00;
              end
              if(_zz_104) begin
                GSHARE_PHT_102 <= 2'b00;
              end
              if(_zz_105) begin
                GSHARE_PHT_103 <= 2'b00;
              end
              if(_zz_106) begin
                GSHARE_PHT_104 <= 2'b00;
              end
              if(_zz_107) begin
                GSHARE_PHT_105 <= 2'b00;
              end
              if(_zz_108) begin
                GSHARE_PHT_106 <= 2'b00;
              end
              if(_zz_109) begin
                GSHARE_PHT_107 <= 2'b00;
              end
              if(_zz_110) begin
                GSHARE_PHT_108 <= 2'b00;
              end
              if(_zz_111) begin
                GSHARE_PHT_109 <= 2'b00;
              end
              if(_zz_112) begin
                GSHARE_PHT_110 <= 2'b00;
              end
              if(_zz_113) begin
                GSHARE_PHT_111 <= 2'b00;
              end
              if(_zz_114) begin
                GSHARE_PHT_112 <= 2'b00;
              end
              if(_zz_115) begin
                GSHARE_PHT_113 <= 2'b00;
              end
              if(_zz_116) begin
                GSHARE_PHT_114 <= 2'b00;
              end
              if(_zz_117) begin
                GSHARE_PHT_115 <= 2'b00;
              end
              if(_zz_118) begin
                GSHARE_PHT_116 <= 2'b00;
              end
              if(_zz_119) begin
                GSHARE_PHT_117 <= 2'b00;
              end
              if(_zz_120) begin
                GSHARE_PHT_118 <= 2'b00;
              end
              if(_zz_121) begin
                GSHARE_PHT_119 <= 2'b00;
              end
              if(_zz_122) begin
                GSHARE_PHT_120 <= 2'b00;
              end
              if(_zz_123) begin
                GSHARE_PHT_121 <= 2'b00;
              end
              if(_zz_124) begin
                GSHARE_PHT_122 <= 2'b00;
              end
              if(_zz_125) begin
                GSHARE_PHT_123 <= 2'b00;
              end
              if(_zz_126) begin
                GSHARE_PHT_124 <= 2'b00;
              end
              if(_zz_127) begin
                GSHARE_PHT_125 <= 2'b00;
              end
              if(_zz_128) begin
                GSHARE_PHT_126 <= 2'b00;
              end
              if(_zz_129) begin
                GSHARE_PHT_127 <= 2'b00;
              end
            end
          end
          2'b10 : begin
            if(train_taken) begin
              if(_zz_2) begin
                GSHARE_PHT_0 <= 2'b11;
              end
              if(_zz_3) begin
                GSHARE_PHT_1 <= 2'b11;
              end
              if(_zz_4) begin
                GSHARE_PHT_2 <= 2'b11;
              end
              if(_zz_5) begin
                GSHARE_PHT_3 <= 2'b11;
              end
              if(_zz_6) begin
                GSHARE_PHT_4 <= 2'b11;
              end
              if(_zz_7) begin
                GSHARE_PHT_5 <= 2'b11;
              end
              if(_zz_8) begin
                GSHARE_PHT_6 <= 2'b11;
              end
              if(_zz_9) begin
                GSHARE_PHT_7 <= 2'b11;
              end
              if(_zz_10) begin
                GSHARE_PHT_8 <= 2'b11;
              end
              if(_zz_11) begin
                GSHARE_PHT_9 <= 2'b11;
              end
              if(_zz_12) begin
                GSHARE_PHT_10 <= 2'b11;
              end
              if(_zz_13) begin
                GSHARE_PHT_11 <= 2'b11;
              end
              if(_zz_14) begin
                GSHARE_PHT_12 <= 2'b11;
              end
              if(_zz_15) begin
                GSHARE_PHT_13 <= 2'b11;
              end
              if(_zz_16) begin
                GSHARE_PHT_14 <= 2'b11;
              end
              if(_zz_17) begin
                GSHARE_PHT_15 <= 2'b11;
              end
              if(_zz_18) begin
                GSHARE_PHT_16 <= 2'b11;
              end
              if(_zz_19) begin
                GSHARE_PHT_17 <= 2'b11;
              end
              if(_zz_20) begin
                GSHARE_PHT_18 <= 2'b11;
              end
              if(_zz_21) begin
                GSHARE_PHT_19 <= 2'b11;
              end
              if(_zz_22) begin
                GSHARE_PHT_20 <= 2'b11;
              end
              if(_zz_23) begin
                GSHARE_PHT_21 <= 2'b11;
              end
              if(_zz_24) begin
                GSHARE_PHT_22 <= 2'b11;
              end
              if(_zz_25) begin
                GSHARE_PHT_23 <= 2'b11;
              end
              if(_zz_26) begin
                GSHARE_PHT_24 <= 2'b11;
              end
              if(_zz_27) begin
                GSHARE_PHT_25 <= 2'b11;
              end
              if(_zz_28) begin
                GSHARE_PHT_26 <= 2'b11;
              end
              if(_zz_29) begin
                GSHARE_PHT_27 <= 2'b11;
              end
              if(_zz_30) begin
                GSHARE_PHT_28 <= 2'b11;
              end
              if(_zz_31) begin
                GSHARE_PHT_29 <= 2'b11;
              end
              if(_zz_32) begin
                GSHARE_PHT_30 <= 2'b11;
              end
              if(_zz_33) begin
                GSHARE_PHT_31 <= 2'b11;
              end
              if(_zz_34) begin
                GSHARE_PHT_32 <= 2'b11;
              end
              if(_zz_35) begin
                GSHARE_PHT_33 <= 2'b11;
              end
              if(_zz_36) begin
                GSHARE_PHT_34 <= 2'b11;
              end
              if(_zz_37) begin
                GSHARE_PHT_35 <= 2'b11;
              end
              if(_zz_38) begin
                GSHARE_PHT_36 <= 2'b11;
              end
              if(_zz_39) begin
                GSHARE_PHT_37 <= 2'b11;
              end
              if(_zz_40) begin
                GSHARE_PHT_38 <= 2'b11;
              end
              if(_zz_41) begin
                GSHARE_PHT_39 <= 2'b11;
              end
              if(_zz_42) begin
                GSHARE_PHT_40 <= 2'b11;
              end
              if(_zz_43) begin
                GSHARE_PHT_41 <= 2'b11;
              end
              if(_zz_44) begin
                GSHARE_PHT_42 <= 2'b11;
              end
              if(_zz_45) begin
                GSHARE_PHT_43 <= 2'b11;
              end
              if(_zz_46) begin
                GSHARE_PHT_44 <= 2'b11;
              end
              if(_zz_47) begin
                GSHARE_PHT_45 <= 2'b11;
              end
              if(_zz_48) begin
                GSHARE_PHT_46 <= 2'b11;
              end
              if(_zz_49) begin
                GSHARE_PHT_47 <= 2'b11;
              end
              if(_zz_50) begin
                GSHARE_PHT_48 <= 2'b11;
              end
              if(_zz_51) begin
                GSHARE_PHT_49 <= 2'b11;
              end
              if(_zz_52) begin
                GSHARE_PHT_50 <= 2'b11;
              end
              if(_zz_53) begin
                GSHARE_PHT_51 <= 2'b11;
              end
              if(_zz_54) begin
                GSHARE_PHT_52 <= 2'b11;
              end
              if(_zz_55) begin
                GSHARE_PHT_53 <= 2'b11;
              end
              if(_zz_56) begin
                GSHARE_PHT_54 <= 2'b11;
              end
              if(_zz_57) begin
                GSHARE_PHT_55 <= 2'b11;
              end
              if(_zz_58) begin
                GSHARE_PHT_56 <= 2'b11;
              end
              if(_zz_59) begin
                GSHARE_PHT_57 <= 2'b11;
              end
              if(_zz_60) begin
                GSHARE_PHT_58 <= 2'b11;
              end
              if(_zz_61) begin
                GSHARE_PHT_59 <= 2'b11;
              end
              if(_zz_62) begin
                GSHARE_PHT_60 <= 2'b11;
              end
              if(_zz_63) begin
                GSHARE_PHT_61 <= 2'b11;
              end
              if(_zz_64) begin
                GSHARE_PHT_62 <= 2'b11;
              end
              if(_zz_65) begin
                GSHARE_PHT_63 <= 2'b11;
              end
              if(_zz_66) begin
                GSHARE_PHT_64 <= 2'b11;
              end
              if(_zz_67) begin
                GSHARE_PHT_65 <= 2'b11;
              end
              if(_zz_68) begin
                GSHARE_PHT_66 <= 2'b11;
              end
              if(_zz_69) begin
                GSHARE_PHT_67 <= 2'b11;
              end
              if(_zz_70) begin
                GSHARE_PHT_68 <= 2'b11;
              end
              if(_zz_71) begin
                GSHARE_PHT_69 <= 2'b11;
              end
              if(_zz_72) begin
                GSHARE_PHT_70 <= 2'b11;
              end
              if(_zz_73) begin
                GSHARE_PHT_71 <= 2'b11;
              end
              if(_zz_74) begin
                GSHARE_PHT_72 <= 2'b11;
              end
              if(_zz_75) begin
                GSHARE_PHT_73 <= 2'b11;
              end
              if(_zz_76) begin
                GSHARE_PHT_74 <= 2'b11;
              end
              if(_zz_77) begin
                GSHARE_PHT_75 <= 2'b11;
              end
              if(_zz_78) begin
                GSHARE_PHT_76 <= 2'b11;
              end
              if(_zz_79) begin
                GSHARE_PHT_77 <= 2'b11;
              end
              if(_zz_80) begin
                GSHARE_PHT_78 <= 2'b11;
              end
              if(_zz_81) begin
                GSHARE_PHT_79 <= 2'b11;
              end
              if(_zz_82) begin
                GSHARE_PHT_80 <= 2'b11;
              end
              if(_zz_83) begin
                GSHARE_PHT_81 <= 2'b11;
              end
              if(_zz_84) begin
                GSHARE_PHT_82 <= 2'b11;
              end
              if(_zz_85) begin
                GSHARE_PHT_83 <= 2'b11;
              end
              if(_zz_86) begin
                GSHARE_PHT_84 <= 2'b11;
              end
              if(_zz_87) begin
                GSHARE_PHT_85 <= 2'b11;
              end
              if(_zz_88) begin
                GSHARE_PHT_86 <= 2'b11;
              end
              if(_zz_89) begin
                GSHARE_PHT_87 <= 2'b11;
              end
              if(_zz_90) begin
                GSHARE_PHT_88 <= 2'b11;
              end
              if(_zz_91) begin
                GSHARE_PHT_89 <= 2'b11;
              end
              if(_zz_92) begin
                GSHARE_PHT_90 <= 2'b11;
              end
              if(_zz_93) begin
                GSHARE_PHT_91 <= 2'b11;
              end
              if(_zz_94) begin
                GSHARE_PHT_92 <= 2'b11;
              end
              if(_zz_95) begin
                GSHARE_PHT_93 <= 2'b11;
              end
              if(_zz_96) begin
                GSHARE_PHT_94 <= 2'b11;
              end
              if(_zz_97) begin
                GSHARE_PHT_95 <= 2'b11;
              end
              if(_zz_98) begin
                GSHARE_PHT_96 <= 2'b11;
              end
              if(_zz_99) begin
                GSHARE_PHT_97 <= 2'b11;
              end
              if(_zz_100) begin
                GSHARE_PHT_98 <= 2'b11;
              end
              if(_zz_101) begin
                GSHARE_PHT_99 <= 2'b11;
              end
              if(_zz_102) begin
                GSHARE_PHT_100 <= 2'b11;
              end
              if(_zz_103) begin
                GSHARE_PHT_101 <= 2'b11;
              end
              if(_zz_104) begin
                GSHARE_PHT_102 <= 2'b11;
              end
              if(_zz_105) begin
                GSHARE_PHT_103 <= 2'b11;
              end
              if(_zz_106) begin
                GSHARE_PHT_104 <= 2'b11;
              end
              if(_zz_107) begin
                GSHARE_PHT_105 <= 2'b11;
              end
              if(_zz_108) begin
                GSHARE_PHT_106 <= 2'b11;
              end
              if(_zz_109) begin
                GSHARE_PHT_107 <= 2'b11;
              end
              if(_zz_110) begin
                GSHARE_PHT_108 <= 2'b11;
              end
              if(_zz_111) begin
                GSHARE_PHT_109 <= 2'b11;
              end
              if(_zz_112) begin
                GSHARE_PHT_110 <= 2'b11;
              end
              if(_zz_113) begin
                GSHARE_PHT_111 <= 2'b11;
              end
              if(_zz_114) begin
                GSHARE_PHT_112 <= 2'b11;
              end
              if(_zz_115) begin
                GSHARE_PHT_113 <= 2'b11;
              end
              if(_zz_116) begin
                GSHARE_PHT_114 <= 2'b11;
              end
              if(_zz_117) begin
                GSHARE_PHT_115 <= 2'b11;
              end
              if(_zz_118) begin
                GSHARE_PHT_116 <= 2'b11;
              end
              if(_zz_119) begin
                GSHARE_PHT_117 <= 2'b11;
              end
              if(_zz_120) begin
                GSHARE_PHT_118 <= 2'b11;
              end
              if(_zz_121) begin
                GSHARE_PHT_119 <= 2'b11;
              end
              if(_zz_122) begin
                GSHARE_PHT_120 <= 2'b11;
              end
              if(_zz_123) begin
                GSHARE_PHT_121 <= 2'b11;
              end
              if(_zz_124) begin
                GSHARE_PHT_122 <= 2'b11;
              end
              if(_zz_125) begin
                GSHARE_PHT_123 <= 2'b11;
              end
              if(_zz_126) begin
                GSHARE_PHT_124 <= 2'b11;
              end
              if(_zz_127) begin
                GSHARE_PHT_125 <= 2'b11;
              end
              if(_zz_128) begin
                GSHARE_PHT_126 <= 2'b11;
              end
              if(_zz_129) begin
                GSHARE_PHT_127 <= 2'b11;
              end
            end else begin
              if(_zz_2) begin
                GSHARE_PHT_0 <= 2'b00;
              end
              if(_zz_3) begin
                GSHARE_PHT_1 <= 2'b00;
              end
              if(_zz_4) begin
                GSHARE_PHT_2 <= 2'b00;
              end
              if(_zz_5) begin
                GSHARE_PHT_3 <= 2'b00;
              end
              if(_zz_6) begin
                GSHARE_PHT_4 <= 2'b00;
              end
              if(_zz_7) begin
                GSHARE_PHT_5 <= 2'b00;
              end
              if(_zz_8) begin
                GSHARE_PHT_6 <= 2'b00;
              end
              if(_zz_9) begin
                GSHARE_PHT_7 <= 2'b00;
              end
              if(_zz_10) begin
                GSHARE_PHT_8 <= 2'b00;
              end
              if(_zz_11) begin
                GSHARE_PHT_9 <= 2'b00;
              end
              if(_zz_12) begin
                GSHARE_PHT_10 <= 2'b00;
              end
              if(_zz_13) begin
                GSHARE_PHT_11 <= 2'b00;
              end
              if(_zz_14) begin
                GSHARE_PHT_12 <= 2'b00;
              end
              if(_zz_15) begin
                GSHARE_PHT_13 <= 2'b00;
              end
              if(_zz_16) begin
                GSHARE_PHT_14 <= 2'b00;
              end
              if(_zz_17) begin
                GSHARE_PHT_15 <= 2'b00;
              end
              if(_zz_18) begin
                GSHARE_PHT_16 <= 2'b00;
              end
              if(_zz_19) begin
                GSHARE_PHT_17 <= 2'b00;
              end
              if(_zz_20) begin
                GSHARE_PHT_18 <= 2'b00;
              end
              if(_zz_21) begin
                GSHARE_PHT_19 <= 2'b00;
              end
              if(_zz_22) begin
                GSHARE_PHT_20 <= 2'b00;
              end
              if(_zz_23) begin
                GSHARE_PHT_21 <= 2'b00;
              end
              if(_zz_24) begin
                GSHARE_PHT_22 <= 2'b00;
              end
              if(_zz_25) begin
                GSHARE_PHT_23 <= 2'b00;
              end
              if(_zz_26) begin
                GSHARE_PHT_24 <= 2'b00;
              end
              if(_zz_27) begin
                GSHARE_PHT_25 <= 2'b00;
              end
              if(_zz_28) begin
                GSHARE_PHT_26 <= 2'b00;
              end
              if(_zz_29) begin
                GSHARE_PHT_27 <= 2'b00;
              end
              if(_zz_30) begin
                GSHARE_PHT_28 <= 2'b00;
              end
              if(_zz_31) begin
                GSHARE_PHT_29 <= 2'b00;
              end
              if(_zz_32) begin
                GSHARE_PHT_30 <= 2'b00;
              end
              if(_zz_33) begin
                GSHARE_PHT_31 <= 2'b00;
              end
              if(_zz_34) begin
                GSHARE_PHT_32 <= 2'b00;
              end
              if(_zz_35) begin
                GSHARE_PHT_33 <= 2'b00;
              end
              if(_zz_36) begin
                GSHARE_PHT_34 <= 2'b00;
              end
              if(_zz_37) begin
                GSHARE_PHT_35 <= 2'b00;
              end
              if(_zz_38) begin
                GSHARE_PHT_36 <= 2'b00;
              end
              if(_zz_39) begin
                GSHARE_PHT_37 <= 2'b00;
              end
              if(_zz_40) begin
                GSHARE_PHT_38 <= 2'b00;
              end
              if(_zz_41) begin
                GSHARE_PHT_39 <= 2'b00;
              end
              if(_zz_42) begin
                GSHARE_PHT_40 <= 2'b00;
              end
              if(_zz_43) begin
                GSHARE_PHT_41 <= 2'b00;
              end
              if(_zz_44) begin
                GSHARE_PHT_42 <= 2'b00;
              end
              if(_zz_45) begin
                GSHARE_PHT_43 <= 2'b00;
              end
              if(_zz_46) begin
                GSHARE_PHT_44 <= 2'b00;
              end
              if(_zz_47) begin
                GSHARE_PHT_45 <= 2'b00;
              end
              if(_zz_48) begin
                GSHARE_PHT_46 <= 2'b00;
              end
              if(_zz_49) begin
                GSHARE_PHT_47 <= 2'b00;
              end
              if(_zz_50) begin
                GSHARE_PHT_48 <= 2'b00;
              end
              if(_zz_51) begin
                GSHARE_PHT_49 <= 2'b00;
              end
              if(_zz_52) begin
                GSHARE_PHT_50 <= 2'b00;
              end
              if(_zz_53) begin
                GSHARE_PHT_51 <= 2'b00;
              end
              if(_zz_54) begin
                GSHARE_PHT_52 <= 2'b00;
              end
              if(_zz_55) begin
                GSHARE_PHT_53 <= 2'b00;
              end
              if(_zz_56) begin
                GSHARE_PHT_54 <= 2'b00;
              end
              if(_zz_57) begin
                GSHARE_PHT_55 <= 2'b00;
              end
              if(_zz_58) begin
                GSHARE_PHT_56 <= 2'b00;
              end
              if(_zz_59) begin
                GSHARE_PHT_57 <= 2'b00;
              end
              if(_zz_60) begin
                GSHARE_PHT_58 <= 2'b00;
              end
              if(_zz_61) begin
                GSHARE_PHT_59 <= 2'b00;
              end
              if(_zz_62) begin
                GSHARE_PHT_60 <= 2'b00;
              end
              if(_zz_63) begin
                GSHARE_PHT_61 <= 2'b00;
              end
              if(_zz_64) begin
                GSHARE_PHT_62 <= 2'b00;
              end
              if(_zz_65) begin
                GSHARE_PHT_63 <= 2'b00;
              end
              if(_zz_66) begin
                GSHARE_PHT_64 <= 2'b00;
              end
              if(_zz_67) begin
                GSHARE_PHT_65 <= 2'b00;
              end
              if(_zz_68) begin
                GSHARE_PHT_66 <= 2'b00;
              end
              if(_zz_69) begin
                GSHARE_PHT_67 <= 2'b00;
              end
              if(_zz_70) begin
                GSHARE_PHT_68 <= 2'b00;
              end
              if(_zz_71) begin
                GSHARE_PHT_69 <= 2'b00;
              end
              if(_zz_72) begin
                GSHARE_PHT_70 <= 2'b00;
              end
              if(_zz_73) begin
                GSHARE_PHT_71 <= 2'b00;
              end
              if(_zz_74) begin
                GSHARE_PHT_72 <= 2'b00;
              end
              if(_zz_75) begin
                GSHARE_PHT_73 <= 2'b00;
              end
              if(_zz_76) begin
                GSHARE_PHT_74 <= 2'b00;
              end
              if(_zz_77) begin
                GSHARE_PHT_75 <= 2'b00;
              end
              if(_zz_78) begin
                GSHARE_PHT_76 <= 2'b00;
              end
              if(_zz_79) begin
                GSHARE_PHT_77 <= 2'b00;
              end
              if(_zz_80) begin
                GSHARE_PHT_78 <= 2'b00;
              end
              if(_zz_81) begin
                GSHARE_PHT_79 <= 2'b00;
              end
              if(_zz_82) begin
                GSHARE_PHT_80 <= 2'b00;
              end
              if(_zz_83) begin
                GSHARE_PHT_81 <= 2'b00;
              end
              if(_zz_84) begin
                GSHARE_PHT_82 <= 2'b00;
              end
              if(_zz_85) begin
                GSHARE_PHT_83 <= 2'b00;
              end
              if(_zz_86) begin
                GSHARE_PHT_84 <= 2'b00;
              end
              if(_zz_87) begin
                GSHARE_PHT_85 <= 2'b00;
              end
              if(_zz_88) begin
                GSHARE_PHT_86 <= 2'b00;
              end
              if(_zz_89) begin
                GSHARE_PHT_87 <= 2'b00;
              end
              if(_zz_90) begin
                GSHARE_PHT_88 <= 2'b00;
              end
              if(_zz_91) begin
                GSHARE_PHT_89 <= 2'b00;
              end
              if(_zz_92) begin
                GSHARE_PHT_90 <= 2'b00;
              end
              if(_zz_93) begin
                GSHARE_PHT_91 <= 2'b00;
              end
              if(_zz_94) begin
                GSHARE_PHT_92 <= 2'b00;
              end
              if(_zz_95) begin
                GSHARE_PHT_93 <= 2'b00;
              end
              if(_zz_96) begin
                GSHARE_PHT_94 <= 2'b00;
              end
              if(_zz_97) begin
                GSHARE_PHT_95 <= 2'b00;
              end
              if(_zz_98) begin
                GSHARE_PHT_96 <= 2'b00;
              end
              if(_zz_99) begin
                GSHARE_PHT_97 <= 2'b00;
              end
              if(_zz_100) begin
                GSHARE_PHT_98 <= 2'b00;
              end
              if(_zz_101) begin
                GSHARE_PHT_99 <= 2'b00;
              end
              if(_zz_102) begin
                GSHARE_PHT_100 <= 2'b00;
              end
              if(_zz_103) begin
                GSHARE_PHT_101 <= 2'b00;
              end
              if(_zz_104) begin
                GSHARE_PHT_102 <= 2'b00;
              end
              if(_zz_105) begin
                GSHARE_PHT_103 <= 2'b00;
              end
              if(_zz_106) begin
                GSHARE_PHT_104 <= 2'b00;
              end
              if(_zz_107) begin
                GSHARE_PHT_105 <= 2'b00;
              end
              if(_zz_108) begin
                GSHARE_PHT_106 <= 2'b00;
              end
              if(_zz_109) begin
                GSHARE_PHT_107 <= 2'b00;
              end
              if(_zz_110) begin
                GSHARE_PHT_108 <= 2'b00;
              end
              if(_zz_111) begin
                GSHARE_PHT_109 <= 2'b00;
              end
              if(_zz_112) begin
                GSHARE_PHT_110 <= 2'b00;
              end
              if(_zz_113) begin
                GSHARE_PHT_111 <= 2'b00;
              end
              if(_zz_114) begin
                GSHARE_PHT_112 <= 2'b00;
              end
              if(_zz_115) begin
                GSHARE_PHT_113 <= 2'b00;
              end
              if(_zz_116) begin
                GSHARE_PHT_114 <= 2'b00;
              end
              if(_zz_117) begin
                GSHARE_PHT_115 <= 2'b00;
              end
              if(_zz_118) begin
                GSHARE_PHT_116 <= 2'b00;
              end
              if(_zz_119) begin
                GSHARE_PHT_117 <= 2'b00;
              end
              if(_zz_120) begin
                GSHARE_PHT_118 <= 2'b00;
              end
              if(_zz_121) begin
                GSHARE_PHT_119 <= 2'b00;
              end
              if(_zz_122) begin
                GSHARE_PHT_120 <= 2'b00;
              end
              if(_zz_123) begin
                GSHARE_PHT_121 <= 2'b00;
              end
              if(_zz_124) begin
                GSHARE_PHT_122 <= 2'b00;
              end
              if(_zz_125) begin
                GSHARE_PHT_123 <= 2'b00;
              end
              if(_zz_126) begin
                GSHARE_PHT_124 <= 2'b00;
              end
              if(_zz_127) begin
                GSHARE_PHT_125 <= 2'b00;
              end
              if(_zz_128) begin
                GSHARE_PHT_126 <= 2'b00;
              end
              if(_zz_129) begin
                GSHARE_PHT_127 <= 2'b00;
              end
            end
          end
          default : begin
            if(when_Predictor_l61) begin
              if(_zz_2) begin
                GSHARE_PHT_0 <= 2'b10;
              end
              if(_zz_3) begin
                GSHARE_PHT_1 <= 2'b10;
              end
              if(_zz_4) begin
                GSHARE_PHT_2 <= 2'b10;
              end
              if(_zz_5) begin
                GSHARE_PHT_3 <= 2'b10;
              end
              if(_zz_6) begin
                GSHARE_PHT_4 <= 2'b10;
              end
              if(_zz_7) begin
                GSHARE_PHT_5 <= 2'b10;
              end
              if(_zz_8) begin
                GSHARE_PHT_6 <= 2'b10;
              end
              if(_zz_9) begin
                GSHARE_PHT_7 <= 2'b10;
              end
              if(_zz_10) begin
                GSHARE_PHT_8 <= 2'b10;
              end
              if(_zz_11) begin
                GSHARE_PHT_9 <= 2'b10;
              end
              if(_zz_12) begin
                GSHARE_PHT_10 <= 2'b10;
              end
              if(_zz_13) begin
                GSHARE_PHT_11 <= 2'b10;
              end
              if(_zz_14) begin
                GSHARE_PHT_12 <= 2'b10;
              end
              if(_zz_15) begin
                GSHARE_PHT_13 <= 2'b10;
              end
              if(_zz_16) begin
                GSHARE_PHT_14 <= 2'b10;
              end
              if(_zz_17) begin
                GSHARE_PHT_15 <= 2'b10;
              end
              if(_zz_18) begin
                GSHARE_PHT_16 <= 2'b10;
              end
              if(_zz_19) begin
                GSHARE_PHT_17 <= 2'b10;
              end
              if(_zz_20) begin
                GSHARE_PHT_18 <= 2'b10;
              end
              if(_zz_21) begin
                GSHARE_PHT_19 <= 2'b10;
              end
              if(_zz_22) begin
                GSHARE_PHT_20 <= 2'b10;
              end
              if(_zz_23) begin
                GSHARE_PHT_21 <= 2'b10;
              end
              if(_zz_24) begin
                GSHARE_PHT_22 <= 2'b10;
              end
              if(_zz_25) begin
                GSHARE_PHT_23 <= 2'b10;
              end
              if(_zz_26) begin
                GSHARE_PHT_24 <= 2'b10;
              end
              if(_zz_27) begin
                GSHARE_PHT_25 <= 2'b10;
              end
              if(_zz_28) begin
                GSHARE_PHT_26 <= 2'b10;
              end
              if(_zz_29) begin
                GSHARE_PHT_27 <= 2'b10;
              end
              if(_zz_30) begin
                GSHARE_PHT_28 <= 2'b10;
              end
              if(_zz_31) begin
                GSHARE_PHT_29 <= 2'b10;
              end
              if(_zz_32) begin
                GSHARE_PHT_30 <= 2'b10;
              end
              if(_zz_33) begin
                GSHARE_PHT_31 <= 2'b10;
              end
              if(_zz_34) begin
                GSHARE_PHT_32 <= 2'b10;
              end
              if(_zz_35) begin
                GSHARE_PHT_33 <= 2'b10;
              end
              if(_zz_36) begin
                GSHARE_PHT_34 <= 2'b10;
              end
              if(_zz_37) begin
                GSHARE_PHT_35 <= 2'b10;
              end
              if(_zz_38) begin
                GSHARE_PHT_36 <= 2'b10;
              end
              if(_zz_39) begin
                GSHARE_PHT_37 <= 2'b10;
              end
              if(_zz_40) begin
                GSHARE_PHT_38 <= 2'b10;
              end
              if(_zz_41) begin
                GSHARE_PHT_39 <= 2'b10;
              end
              if(_zz_42) begin
                GSHARE_PHT_40 <= 2'b10;
              end
              if(_zz_43) begin
                GSHARE_PHT_41 <= 2'b10;
              end
              if(_zz_44) begin
                GSHARE_PHT_42 <= 2'b10;
              end
              if(_zz_45) begin
                GSHARE_PHT_43 <= 2'b10;
              end
              if(_zz_46) begin
                GSHARE_PHT_44 <= 2'b10;
              end
              if(_zz_47) begin
                GSHARE_PHT_45 <= 2'b10;
              end
              if(_zz_48) begin
                GSHARE_PHT_46 <= 2'b10;
              end
              if(_zz_49) begin
                GSHARE_PHT_47 <= 2'b10;
              end
              if(_zz_50) begin
                GSHARE_PHT_48 <= 2'b10;
              end
              if(_zz_51) begin
                GSHARE_PHT_49 <= 2'b10;
              end
              if(_zz_52) begin
                GSHARE_PHT_50 <= 2'b10;
              end
              if(_zz_53) begin
                GSHARE_PHT_51 <= 2'b10;
              end
              if(_zz_54) begin
                GSHARE_PHT_52 <= 2'b10;
              end
              if(_zz_55) begin
                GSHARE_PHT_53 <= 2'b10;
              end
              if(_zz_56) begin
                GSHARE_PHT_54 <= 2'b10;
              end
              if(_zz_57) begin
                GSHARE_PHT_55 <= 2'b10;
              end
              if(_zz_58) begin
                GSHARE_PHT_56 <= 2'b10;
              end
              if(_zz_59) begin
                GSHARE_PHT_57 <= 2'b10;
              end
              if(_zz_60) begin
                GSHARE_PHT_58 <= 2'b10;
              end
              if(_zz_61) begin
                GSHARE_PHT_59 <= 2'b10;
              end
              if(_zz_62) begin
                GSHARE_PHT_60 <= 2'b10;
              end
              if(_zz_63) begin
                GSHARE_PHT_61 <= 2'b10;
              end
              if(_zz_64) begin
                GSHARE_PHT_62 <= 2'b10;
              end
              if(_zz_65) begin
                GSHARE_PHT_63 <= 2'b10;
              end
              if(_zz_66) begin
                GSHARE_PHT_64 <= 2'b10;
              end
              if(_zz_67) begin
                GSHARE_PHT_65 <= 2'b10;
              end
              if(_zz_68) begin
                GSHARE_PHT_66 <= 2'b10;
              end
              if(_zz_69) begin
                GSHARE_PHT_67 <= 2'b10;
              end
              if(_zz_70) begin
                GSHARE_PHT_68 <= 2'b10;
              end
              if(_zz_71) begin
                GSHARE_PHT_69 <= 2'b10;
              end
              if(_zz_72) begin
                GSHARE_PHT_70 <= 2'b10;
              end
              if(_zz_73) begin
                GSHARE_PHT_71 <= 2'b10;
              end
              if(_zz_74) begin
                GSHARE_PHT_72 <= 2'b10;
              end
              if(_zz_75) begin
                GSHARE_PHT_73 <= 2'b10;
              end
              if(_zz_76) begin
                GSHARE_PHT_74 <= 2'b10;
              end
              if(_zz_77) begin
                GSHARE_PHT_75 <= 2'b10;
              end
              if(_zz_78) begin
                GSHARE_PHT_76 <= 2'b10;
              end
              if(_zz_79) begin
                GSHARE_PHT_77 <= 2'b10;
              end
              if(_zz_80) begin
                GSHARE_PHT_78 <= 2'b10;
              end
              if(_zz_81) begin
                GSHARE_PHT_79 <= 2'b10;
              end
              if(_zz_82) begin
                GSHARE_PHT_80 <= 2'b10;
              end
              if(_zz_83) begin
                GSHARE_PHT_81 <= 2'b10;
              end
              if(_zz_84) begin
                GSHARE_PHT_82 <= 2'b10;
              end
              if(_zz_85) begin
                GSHARE_PHT_83 <= 2'b10;
              end
              if(_zz_86) begin
                GSHARE_PHT_84 <= 2'b10;
              end
              if(_zz_87) begin
                GSHARE_PHT_85 <= 2'b10;
              end
              if(_zz_88) begin
                GSHARE_PHT_86 <= 2'b10;
              end
              if(_zz_89) begin
                GSHARE_PHT_87 <= 2'b10;
              end
              if(_zz_90) begin
                GSHARE_PHT_88 <= 2'b10;
              end
              if(_zz_91) begin
                GSHARE_PHT_89 <= 2'b10;
              end
              if(_zz_92) begin
                GSHARE_PHT_90 <= 2'b10;
              end
              if(_zz_93) begin
                GSHARE_PHT_91 <= 2'b10;
              end
              if(_zz_94) begin
                GSHARE_PHT_92 <= 2'b10;
              end
              if(_zz_95) begin
                GSHARE_PHT_93 <= 2'b10;
              end
              if(_zz_96) begin
                GSHARE_PHT_94 <= 2'b10;
              end
              if(_zz_97) begin
                GSHARE_PHT_95 <= 2'b10;
              end
              if(_zz_98) begin
                GSHARE_PHT_96 <= 2'b10;
              end
              if(_zz_99) begin
                GSHARE_PHT_97 <= 2'b10;
              end
              if(_zz_100) begin
                GSHARE_PHT_98 <= 2'b10;
              end
              if(_zz_101) begin
                GSHARE_PHT_99 <= 2'b10;
              end
              if(_zz_102) begin
                GSHARE_PHT_100 <= 2'b10;
              end
              if(_zz_103) begin
                GSHARE_PHT_101 <= 2'b10;
              end
              if(_zz_104) begin
                GSHARE_PHT_102 <= 2'b10;
              end
              if(_zz_105) begin
                GSHARE_PHT_103 <= 2'b10;
              end
              if(_zz_106) begin
                GSHARE_PHT_104 <= 2'b10;
              end
              if(_zz_107) begin
                GSHARE_PHT_105 <= 2'b10;
              end
              if(_zz_108) begin
                GSHARE_PHT_106 <= 2'b10;
              end
              if(_zz_109) begin
                GSHARE_PHT_107 <= 2'b10;
              end
              if(_zz_110) begin
                GSHARE_PHT_108 <= 2'b10;
              end
              if(_zz_111) begin
                GSHARE_PHT_109 <= 2'b10;
              end
              if(_zz_112) begin
                GSHARE_PHT_110 <= 2'b10;
              end
              if(_zz_113) begin
                GSHARE_PHT_111 <= 2'b10;
              end
              if(_zz_114) begin
                GSHARE_PHT_112 <= 2'b10;
              end
              if(_zz_115) begin
                GSHARE_PHT_113 <= 2'b10;
              end
              if(_zz_116) begin
                GSHARE_PHT_114 <= 2'b10;
              end
              if(_zz_117) begin
                GSHARE_PHT_115 <= 2'b10;
              end
              if(_zz_118) begin
                GSHARE_PHT_116 <= 2'b10;
              end
              if(_zz_119) begin
                GSHARE_PHT_117 <= 2'b10;
              end
              if(_zz_120) begin
                GSHARE_PHT_118 <= 2'b10;
              end
              if(_zz_121) begin
                GSHARE_PHT_119 <= 2'b10;
              end
              if(_zz_122) begin
                GSHARE_PHT_120 <= 2'b10;
              end
              if(_zz_123) begin
                GSHARE_PHT_121 <= 2'b10;
              end
              if(_zz_124) begin
                GSHARE_PHT_122 <= 2'b10;
              end
              if(_zz_125) begin
                GSHARE_PHT_123 <= 2'b10;
              end
              if(_zz_126) begin
                GSHARE_PHT_124 <= 2'b10;
              end
              if(_zz_127) begin
                GSHARE_PHT_125 <= 2'b10;
              end
              if(_zz_128) begin
                GSHARE_PHT_126 <= 2'b10;
              end
              if(_zz_129) begin
                GSHARE_PHT_127 <= 2'b10;
              end
            end else begin
              if(_zz_2) begin
                GSHARE_PHT_0 <= 2'b11;
              end
              if(_zz_3) begin
                GSHARE_PHT_1 <= 2'b11;
              end
              if(_zz_4) begin
                GSHARE_PHT_2 <= 2'b11;
              end
              if(_zz_5) begin
                GSHARE_PHT_3 <= 2'b11;
              end
              if(_zz_6) begin
                GSHARE_PHT_4 <= 2'b11;
              end
              if(_zz_7) begin
                GSHARE_PHT_5 <= 2'b11;
              end
              if(_zz_8) begin
                GSHARE_PHT_6 <= 2'b11;
              end
              if(_zz_9) begin
                GSHARE_PHT_7 <= 2'b11;
              end
              if(_zz_10) begin
                GSHARE_PHT_8 <= 2'b11;
              end
              if(_zz_11) begin
                GSHARE_PHT_9 <= 2'b11;
              end
              if(_zz_12) begin
                GSHARE_PHT_10 <= 2'b11;
              end
              if(_zz_13) begin
                GSHARE_PHT_11 <= 2'b11;
              end
              if(_zz_14) begin
                GSHARE_PHT_12 <= 2'b11;
              end
              if(_zz_15) begin
                GSHARE_PHT_13 <= 2'b11;
              end
              if(_zz_16) begin
                GSHARE_PHT_14 <= 2'b11;
              end
              if(_zz_17) begin
                GSHARE_PHT_15 <= 2'b11;
              end
              if(_zz_18) begin
                GSHARE_PHT_16 <= 2'b11;
              end
              if(_zz_19) begin
                GSHARE_PHT_17 <= 2'b11;
              end
              if(_zz_20) begin
                GSHARE_PHT_18 <= 2'b11;
              end
              if(_zz_21) begin
                GSHARE_PHT_19 <= 2'b11;
              end
              if(_zz_22) begin
                GSHARE_PHT_20 <= 2'b11;
              end
              if(_zz_23) begin
                GSHARE_PHT_21 <= 2'b11;
              end
              if(_zz_24) begin
                GSHARE_PHT_22 <= 2'b11;
              end
              if(_zz_25) begin
                GSHARE_PHT_23 <= 2'b11;
              end
              if(_zz_26) begin
                GSHARE_PHT_24 <= 2'b11;
              end
              if(_zz_27) begin
                GSHARE_PHT_25 <= 2'b11;
              end
              if(_zz_28) begin
                GSHARE_PHT_26 <= 2'b11;
              end
              if(_zz_29) begin
                GSHARE_PHT_27 <= 2'b11;
              end
              if(_zz_30) begin
                GSHARE_PHT_28 <= 2'b11;
              end
              if(_zz_31) begin
                GSHARE_PHT_29 <= 2'b11;
              end
              if(_zz_32) begin
                GSHARE_PHT_30 <= 2'b11;
              end
              if(_zz_33) begin
                GSHARE_PHT_31 <= 2'b11;
              end
              if(_zz_34) begin
                GSHARE_PHT_32 <= 2'b11;
              end
              if(_zz_35) begin
                GSHARE_PHT_33 <= 2'b11;
              end
              if(_zz_36) begin
                GSHARE_PHT_34 <= 2'b11;
              end
              if(_zz_37) begin
                GSHARE_PHT_35 <= 2'b11;
              end
              if(_zz_38) begin
                GSHARE_PHT_36 <= 2'b11;
              end
              if(_zz_39) begin
                GSHARE_PHT_37 <= 2'b11;
              end
              if(_zz_40) begin
                GSHARE_PHT_38 <= 2'b11;
              end
              if(_zz_41) begin
                GSHARE_PHT_39 <= 2'b11;
              end
              if(_zz_42) begin
                GSHARE_PHT_40 <= 2'b11;
              end
              if(_zz_43) begin
                GSHARE_PHT_41 <= 2'b11;
              end
              if(_zz_44) begin
                GSHARE_PHT_42 <= 2'b11;
              end
              if(_zz_45) begin
                GSHARE_PHT_43 <= 2'b11;
              end
              if(_zz_46) begin
                GSHARE_PHT_44 <= 2'b11;
              end
              if(_zz_47) begin
                GSHARE_PHT_45 <= 2'b11;
              end
              if(_zz_48) begin
                GSHARE_PHT_46 <= 2'b11;
              end
              if(_zz_49) begin
                GSHARE_PHT_47 <= 2'b11;
              end
              if(_zz_50) begin
                GSHARE_PHT_48 <= 2'b11;
              end
              if(_zz_51) begin
                GSHARE_PHT_49 <= 2'b11;
              end
              if(_zz_52) begin
                GSHARE_PHT_50 <= 2'b11;
              end
              if(_zz_53) begin
                GSHARE_PHT_51 <= 2'b11;
              end
              if(_zz_54) begin
                GSHARE_PHT_52 <= 2'b11;
              end
              if(_zz_55) begin
                GSHARE_PHT_53 <= 2'b11;
              end
              if(_zz_56) begin
                GSHARE_PHT_54 <= 2'b11;
              end
              if(_zz_57) begin
                GSHARE_PHT_55 <= 2'b11;
              end
              if(_zz_58) begin
                GSHARE_PHT_56 <= 2'b11;
              end
              if(_zz_59) begin
                GSHARE_PHT_57 <= 2'b11;
              end
              if(_zz_60) begin
                GSHARE_PHT_58 <= 2'b11;
              end
              if(_zz_61) begin
                GSHARE_PHT_59 <= 2'b11;
              end
              if(_zz_62) begin
                GSHARE_PHT_60 <= 2'b11;
              end
              if(_zz_63) begin
                GSHARE_PHT_61 <= 2'b11;
              end
              if(_zz_64) begin
                GSHARE_PHT_62 <= 2'b11;
              end
              if(_zz_65) begin
                GSHARE_PHT_63 <= 2'b11;
              end
              if(_zz_66) begin
                GSHARE_PHT_64 <= 2'b11;
              end
              if(_zz_67) begin
                GSHARE_PHT_65 <= 2'b11;
              end
              if(_zz_68) begin
                GSHARE_PHT_66 <= 2'b11;
              end
              if(_zz_69) begin
                GSHARE_PHT_67 <= 2'b11;
              end
              if(_zz_70) begin
                GSHARE_PHT_68 <= 2'b11;
              end
              if(_zz_71) begin
                GSHARE_PHT_69 <= 2'b11;
              end
              if(_zz_72) begin
                GSHARE_PHT_70 <= 2'b11;
              end
              if(_zz_73) begin
                GSHARE_PHT_71 <= 2'b11;
              end
              if(_zz_74) begin
                GSHARE_PHT_72 <= 2'b11;
              end
              if(_zz_75) begin
                GSHARE_PHT_73 <= 2'b11;
              end
              if(_zz_76) begin
                GSHARE_PHT_74 <= 2'b11;
              end
              if(_zz_77) begin
                GSHARE_PHT_75 <= 2'b11;
              end
              if(_zz_78) begin
                GSHARE_PHT_76 <= 2'b11;
              end
              if(_zz_79) begin
                GSHARE_PHT_77 <= 2'b11;
              end
              if(_zz_80) begin
                GSHARE_PHT_78 <= 2'b11;
              end
              if(_zz_81) begin
                GSHARE_PHT_79 <= 2'b11;
              end
              if(_zz_82) begin
                GSHARE_PHT_80 <= 2'b11;
              end
              if(_zz_83) begin
                GSHARE_PHT_81 <= 2'b11;
              end
              if(_zz_84) begin
                GSHARE_PHT_82 <= 2'b11;
              end
              if(_zz_85) begin
                GSHARE_PHT_83 <= 2'b11;
              end
              if(_zz_86) begin
                GSHARE_PHT_84 <= 2'b11;
              end
              if(_zz_87) begin
                GSHARE_PHT_85 <= 2'b11;
              end
              if(_zz_88) begin
                GSHARE_PHT_86 <= 2'b11;
              end
              if(_zz_89) begin
                GSHARE_PHT_87 <= 2'b11;
              end
              if(_zz_90) begin
                GSHARE_PHT_88 <= 2'b11;
              end
              if(_zz_91) begin
                GSHARE_PHT_89 <= 2'b11;
              end
              if(_zz_92) begin
                GSHARE_PHT_90 <= 2'b11;
              end
              if(_zz_93) begin
                GSHARE_PHT_91 <= 2'b11;
              end
              if(_zz_94) begin
                GSHARE_PHT_92 <= 2'b11;
              end
              if(_zz_95) begin
                GSHARE_PHT_93 <= 2'b11;
              end
              if(_zz_96) begin
                GSHARE_PHT_94 <= 2'b11;
              end
              if(_zz_97) begin
                GSHARE_PHT_95 <= 2'b11;
              end
              if(_zz_98) begin
                GSHARE_PHT_96 <= 2'b11;
              end
              if(_zz_99) begin
                GSHARE_PHT_97 <= 2'b11;
              end
              if(_zz_100) begin
                GSHARE_PHT_98 <= 2'b11;
              end
              if(_zz_101) begin
                GSHARE_PHT_99 <= 2'b11;
              end
              if(_zz_102) begin
                GSHARE_PHT_100 <= 2'b11;
              end
              if(_zz_103) begin
                GSHARE_PHT_101 <= 2'b11;
              end
              if(_zz_104) begin
                GSHARE_PHT_102 <= 2'b11;
              end
              if(_zz_105) begin
                GSHARE_PHT_103 <= 2'b11;
              end
              if(_zz_106) begin
                GSHARE_PHT_104 <= 2'b11;
              end
              if(_zz_107) begin
                GSHARE_PHT_105 <= 2'b11;
              end
              if(_zz_108) begin
                GSHARE_PHT_106 <= 2'b11;
              end
              if(_zz_109) begin
                GSHARE_PHT_107 <= 2'b11;
              end
              if(_zz_110) begin
                GSHARE_PHT_108 <= 2'b11;
              end
              if(_zz_111) begin
                GSHARE_PHT_109 <= 2'b11;
              end
              if(_zz_112) begin
                GSHARE_PHT_110 <= 2'b11;
              end
              if(_zz_113) begin
                GSHARE_PHT_111 <= 2'b11;
              end
              if(_zz_114) begin
                GSHARE_PHT_112 <= 2'b11;
              end
              if(_zz_115) begin
                GSHARE_PHT_113 <= 2'b11;
              end
              if(_zz_116) begin
                GSHARE_PHT_114 <= 2'b11;
              end
              if(_zz_117) begin
                GSHARE_PHT_115 <= 2'b11;
              end
              if(_zz_118) begin
                GSHARE_PHT_116 <= 2'b11;
              end
              if(_zz_119) begin
                GSHARE_PHT_117 <= 2'b11;
              end
              if(_zz_120) begin
                GSHARE_PHT_118 <= 2'b11;
              end
              if(_zz_121) begin
                GSHARE_PHT_119 <= 2'b11;
              end
              if(_zz_122) begin
                GSHARE_PHT_120 <= 2'b11;
              end
              if(_zz_123) begin
                GSHARE_PHT_121 <= 2'b11;
              end
              if(_zz_124) begin
                GSHARE_PHT_122 <= 2'b11;
              end
              if(_zz_125) begin
                GSHARE_PHT_123 <= 2'b11;
              end
              if(_zz_126) begin
                GSHARE_PHT_124 <= 2'b11;
              end
              if(_zz_127) begin
                GSHARE_PHT_125 <= 2'b11;
              end
              if(_zz_128) begin
                GSHARE_PHT_126 <= 2'b11;
              end
              if(_zz_129) begin
                GSHARE_PHT_127 <= 2'b11;
              end
            end
          end
        endcase
      end
      if(when_Predictor_l70) begin
        GSHARE_global_branch_history <= {train_history[5 : 0],train_taken};
      end else begin
        if(predict_valid) begin
          GSHARE_global_branch_history <= {GSHARE_global_branch_history[5 : 0],predict_taken};
        end
      end
      BTB_btb_alloc_index_value <= BTB_btb_alloc_index_valueNext;
      if(BTB_btb_is_hit) begin
        if(_zz_130[0]) begin
          BTB_source_pc_0 <= train_pc;
        end
        if(_zz_130[1]) begin
          BTB_source_pc_1 <= train_pc;
        end
        if(_zz_130[2]) begin
          BTB_source_pc_2 <= train_pc;
        end
        if(_zz_130[3]) begin
          BTB_source_pc_3 <= train_pc;
        end
        BTB_call[BTB_btb_write_index] <= train_is_call;
        BTB_ret[BTB_btb_write_index] <= train_is_ret;
        BTB_jmp[BTB_btb_write_index] <= train_is_jmp;
        if(_zz_131[0]) begin
          BTB_target_pc_0 <= train_pc_next;
        end
        if(_zz_131[1]) begin
          BTB_target_pc_1 <= train_pc_next;
        end
        if(_zz_131[2]) begin
          BTB_target_pc_2 <= train_pc_next;
        end
        if(_zz_131[3]) begin
          BTB_target_pc_3 <= train_pc_next;
        end
      end else begin
        if(BTB_btb_is_miss) begin
          BTB_valid[BTB_btb_alloc_index_value] <= 1'b1;
          if(_zz_132[0]) begin
            BTB_source_pc_0 <= train_pc;
          end
          if(_zz_132[1]) begin
            BTB_source_pc_1 <= train_pc;
          end
          if(_zz_132[2]) begin
            BTB_source_pc_2 <= train_pc;
          end
          if(_zz_132[3]) begin
            BTB_source_pc_3 <= train_pc;
          end
          BTB_call[BTB_btb_alloc_index_value] <= train_is_call;
          BTB_ret[BTB_btb_alloc_index_value] <= train_is_ret;
          BTB_jmp[BTB_btb_alloc_index_value] <= train_is_jmp;
          if(_zz_133[0]) begin
            BTB_target_pc_0 <= train_pc_next;
          end
          if(_zz_133[1]) begin
            BTB_target_pc_1 <= train_pc_next;
          end
          if(_zz_133[2]) begin
            BTB_target_pc_2 <= train_pc_next;
          end
          if(_zz_133[3]) begin
            BTB_target_pc_3 <= train_pc_next;
          end
        end
      end
      RAS_ras_curr_index_proven <= RAS_ras_next_index;
      if(when_Predictor_l197) begin
        RAS_ras_curr_index <= RAS_ras_next_index;
      end else begin
        if(RAS_ras_call_matched) begin
          RAS_ras_curr_index <= RAS_ras_next_index;
        end else begin
          if(when_Predictor_l205) begin
            RAS_ras_curr_index <= RAS_ras_next_index;
          end else begin
            if(RAS_ras_ret_matched) begin
              RAS_ras_curr_index <= RAS_ras_next_index;
            end
          end
        end
      end
    end
  end

  always @(posedge clk) begin
    if(when_Predictor_l197) begin
      if(_zz_135) begin
        RAS_ras_regfile_0 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_136) begin
        RAS_ras_regfile_1 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_137) begin
        RAS_ras_regfile_2 <= _zz_RAS_ras_regfile_0;
      end
      if(_zz_138) begin
        RAS_ras_regfile_3 <= _zz_RAS_ras_regfile_0;
      end
    end else begin
      if(RAS_ras_call_matched) begin
        if(_zz_135) begin
          RAS_ras_regfile_0 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_136) begin
          RAS_ras_regfile_1 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_137) begin
          RAS_ras_regfile_2 <= _zz_RAS_ras_regfile_0_1;
        end
        if(_zz_138) begin
          RAS_ras_regfile_3 <= _zz_RAS_ras_regfile_0_1;
        end
      end
    end
  end


endmodule

module FIFO_2 (
  input               ports_s_ports_valid,
  output              ports_s_ports_ready,
  input      [31:0]   ports_s_ports_payload,
  output              ports_m_ports_valid,
  input               ports_m_ports_ready,
  output     [31:0]   ports_m_ports_payload,
  input               flush,
  input               clk,
  input               reset
);

  reg        [31:0]   _zz_ports_m_ports_payload;
  reg        [2:0]    read_ptr;
  reg        [2:0]    write_ptr;
  wire       [1:0]    read_addr;
  wire       [1:0]    next_read_addr;
  wire       [1:0]    write_addr;
  wire                fifo_empty;
  wire                fifo_full;
  reg        [31:0]   fifo_ram_0;
  reg        [31:0]   fifo_ram_1;
  reg        [31:0]   fifo_ram_2;
  reg        [31:0]   fifo_ram_3;
  wire                ports_m_ports_fire;
  wire       [3:0]    _zz_1;
  wire                ports_s_ports_fire;

  always @(*) begin
    case(read_addr)
      2'b00 : _zz_ports_m_ports_payload = fifo_ram_0;
      2'b01 : _zz_ports_m_ports_payload = fifo_ram_1;
      2'b10 : _zz_ports_m_ports_payload = fifo_ram_2;
      default : _zz_ports_m_ports_payload = fifo_ram_3;
    endcase
  end

  assign read_addr = read_ptr[1 : 0];
  assign next_read_addr = (read_addr + 2'b01);
  assign write_addr = write_ptr[1 : 0];
  assign fifo_empty = (read_ptr == write_ptr);
  assign fifo_full = ((read_addr == write_addr) && (read_ptr[2] != write_ptr[2]));
  assign ports_m_ports_fire = (ports_m_ports_valid && ports_m_ports_ready);
  assign _zz_1 = ({3'd0,1'b1} <<< write_addr);
  assign ports_s_ports_fire = (ports_s_ports_valid && ports_s_ports_ready);
  assign ports_s_ports_ready = (! fifo_full);
  assign ports_m_ports_valid = (! fifo_empty);
  assign ports_m_ports_payload = _zz_ports_m_ports_payload;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      read_ptr <= 3'b000;
      write_ptr <= 3'b000;
    end else begin
      if(flush) begin
        read_ptr <= 3'b000;
      end else begin
        if(ports_m_ports_fire) begin
          read_ptr <= (read_ptr + 3'b001);
        end
      end
      if(flush) begin
        write_ptr <= 3'b000;
      end else begin
        if(ports_s_ports_fire) begin
          write_ptr <= (write_ptr + 3'b001);
        end
      end
    end
  end

  always @(posedge clk) begin
    if(!flush) begin
      if(ports_s_ports_fire) begin
        if(_zz_1[0]) begin
          fifo_ram_0 <= ports_s_ports_payload;
        end
        if(_zz_1[1]) begin
          fifo_ram_1 <= ports_s_ports_payload;
        end
        if(_zz_1[2]) begin
          fifo_ram_2 <= ports_s_ports_payload;
        end
        if(_zz_1[3]) begin
          fifo_ram_3 <= ports_s_ports_payload;
        end
      end
    end
  end


endmodule

module FIFO_1 (
  input               ports_s_ports_valid,
  output              ports_s_ports_ready,
  input               ports_s_ports_payload,
  output              ports_m_ports_valid,
  input               ports_m_ports_ready,
  output              ports_m_ports_payload,
  input               flush,
  input               clk,
  input               reset
);

  reg                 _zz_ports_m_ports_payload;
  reg        [2:0]    read_ptr;
  reg        [2:0]    write_ptr;
  wire       [1:0]    read_addr;
  wire       [1:0]    next_read_addr;
  wire       [1:0]    write_addr;
  wire                fifo_empty;
  wire                fifo_full;
  reg                 fifo_ram_0;
  reg                 fifo_ram_1;
  reg                 fifo_ram_2;
  reg                 fifo_ram_3;
  wire                ports_m_ports_fire;
  wire       [3:0]    _zz_1;
  wire                ports_s_ports_fire;

  always @(*) begin
    case(read_addr)
      2'b00 : _zz_ports_m_ports_payload = fifo_ram_0;
      2'b01 : _zz_ports_m_ports_payload = fifo_ram_1;
      2'b10 : _zz_ports_m_ports_payload = fifo_ram_2;
      default : _zz_ports_m_ports_payload = fifo_ram_3;
    endcase
  end

  assign read_addr = read_ptr[1 : 0];
  assign next_read_addr = (read_addr + 2'b01);
  assign write_addr = write_ptr[1 : 0];
  assign fifo_empty = (read_ptr == write_ptr);
  assign fifo_full = ((read_addr == write_addr) && (read_ptr[2] != write_ptr[2]));
  assign ports_m_ports_fire = (ports_m_ports_valid && ports_m_ports_ready);
  assign _zz_1 = ({3'd0,1'b1} <<< write_addr);
  assign ports_s_ports_fire = (ports_s_ports_valid && ports_s_ports_ready);
  assign ports_s_ports_ready = (! fifo_full);
  assign ports_m_ports_valid = (! fifo_empty);
  assign ports_m_ports_payload = _zz_ports_m_ports_payload;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      read_ptr <= 3'b000;
      write_ptr <= 3'b000;
    end else begin
      if(flush) begin
        read_ptr <= 3'b000;
      end else begin
        if(ports_m_ports_fire) begin
          read_ptr <= (read_ptr + 3'b001);
        end
      end
      if(flush) begin
        write_ptr <= 3'b000;
      end else begin
        if(ports_s_ports_fire) begin
          write_ptr <= (write_ptr + 3'b001);
        end
      end
    end
  end

  always @(posedge clk) begin
    if(!flush) begin
      if(ports_s_ports_fire) begin
        if(_zz_1[0]) begin
          fifo_ram_0 <= ports_s_ports_payload;
        end
        if(_zz_1[1]) begin
          fifo_ram_1 <= ports_s_ports_payload;
        end
        if(_zz_1[2]) begin
          fifo_ram_2 <= ports_s_ports_payload;
        end
        if(_zz_1[3]) begin
          fifo_ram_3 <= ports_s_ports_payload;
        end
      end
    end
  end


endmodule

module FIFO (
  input               ports_s_ports_valid,
  output              ports_s_ports_ready,
  input      [63:0]   ports_s_ports_payload,
  output              ports_m_ports_valid,
  input               ports_m_ports_ready,
  output     [63:0]   ports_m_ports_payload,
  input               flush,
  output     [63:0]   next_payload,
  output              next_valid,
  input               clk,
  input               reset
);

  reg        [63:0]   _zz_ports_m_ports_payload;
  reg        [63:0]   _zz_next_payload;
  reg        [2:0]    read_ptr;
  reg        [2:0]    write_ptr;
  wire       [1:0]    read_addr;
  wire       [1:0]    next_read_addr;
  wire       [1:0]    write_addr;
  wire                fifo_empty;
  wire                fifo_full;
  reg        [63:0]   fifo_ram_0;
  reg        [63:0]   fifo_ram_1;
  reg        [63:0]   fifo_ram_2;
  reg        [63:0]   fifo_ram_3;
  wire                ports_m_ports_fire;
  wire       [3:0]    _zz_1;
  wire                ports_s_ports_fire;
  reg        [2:0]    fifo_cnt;
  wire                ports_s_ports_fire_1;
  wire                ports_m_ports_fire_1;
  wire                when_FIFO_l61;
  wire                ports_s_ports_fire_2;
  wire                ports_m_ports_fire_2;
  wire                when_FIFO_l64;

  always @(*) begin
    case(read_addr)
      2'b00 : _zz_ports_m_ports_payload = fifo_ram_0;
      2'b01 : _zz_ports_m_ports_payload = fifo_ram_1;
      2'b10 : _zz_ports_m_ports_payload = fifo_ram_2;
      default : _zz_ports_m_ports_payload = fifo_ram_3;
    endcase
  end

  always @(*) begin
    case(next_read_addr)
      2'b00 : _zz_next_payload = fifo_ram_0;
      2'b01 : _zz_next_payload = fifo_ram_1;
      2'b10 : _zz_next_payload = fifo_ram_2;
      default : _zz_next_payload = fifo_ram_3;
    endcase
  end

  assign read_addr = read_ptr[1 : 0];
  assign next_read_addr = (read_addr + 2'b01);
  assign write_addr = write_ptr[1 : 0];
  assign fifo_empty = (read_ptr == write_ptr);
  assign fifo_full = ((read_addr == write_addr) && (read_ptr[2] != write_ptr[2]));
  assign ports_m_ports_fire = (ports_m_ports_valid && ports_m_ports_ready);
  assign _zz_1 = ({3'd0,1'b1} <<< write_addr);
  assign ports_s_ports_fire = (ports_s_ports_valid && ports_s_ports_ready);
  assign ports_s_ports_ready = (! fifo_full);
  assign ports_m_ports_valid = (! fifo_empty);
  assign ports_m_ports_payload = _zz_ports_m_ports_payload;
  assign next_payload = _zz_next_payload;
  assign ports_s_ports_fire_1 = (ports_s_ports_valid && ports_s_ports_ready);
  assign ports_m_ports_fire_1 = (ports_m_ports_valid && ports_m_ports_ready);
  assign when_FIFO_l61 = (ports_s_ports_fire_1 && (! ports_m_ports_fire_1));
  assign ports_s_ports_fire_2 = (ports_s_ports_valid && ports_s_ports_ready);
  assign ports_m_ports_fire_2 = (ports_m_ports_valid && ports_m_ports_ready);
  assign when_FIFO_l64 = ((! ports_s_ports_fire_2) && ports_m_ports_fire_2);
  assign next_valid = (3'b010 <= fifo_cnt);
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      read_ptr <= 3'b000;
      write_ptr <= 3'b000;
      fifo_cnt <= 3'b000;
    end else begin
      if(flush) begin
        read_ptr <= 3'b000;
      end else begin
        if(ports_m_ports_fire) begin
          read_ptr <= (read_ptr + 3'b001);
        end
      end
      if(flush) begin
        write_ptr <= 3'b000;
      end else begin
        if(ports_s_ports_fire) begin
          write_ptr <= (write_ptr + 3'b001);
        end
      end
      if(flush) begin
        fifo_cnt <= 3'b000;
      end else begin
        if(when_FIFO_l61) begin
          fifo_cnt <= (fifo_cnt + 3'b001);
        end else begin
          if(when_FIFO_l64) begin
            fifo_cnt <= (fifo_cnt - 3'b001);
          end
        end
      end
    end
  end

  always @(posedge clk) begin
    if(!flush) begin
      if(ports_s_ports_fire) begin
        if(_zz_1[0]) begin
          fifo_ram_0 <= ports_s_ports_payload;
        end
        if(_zz_1[1]) begin
          fifo_ram_1 <= ports_s_ports_payload;
        end
        if(_zz_1[2]) begin
          fifo_ram_2 <= ports_s_ports_payload;
        end
        if(_zz_1[3]) begin
          fifo_ram_3 <= ports_s_ports_payload;
        end
      end
    end
  end


endmodule
